module mvt_float(
	input clk,
	input rst,

	input [0 : 0]start_in,
	input start_valid,
	output start_ready,

	output [0 : 0]end_out,
	output end_valid,
	input end_ready,

	output [5 : 0]x1_address0,
	output x1_ce0,
	output x1_we0,
	output [31 : 0]x1_dout0,
	input [31 : 0]x1_din0,
	output [5 : 0]x1_address1,
	output x1_ce1,
	output x1_we1,
	output [31 : 0]x1_dout1,
	input [31 : 0]x1_din1,

	output [11 : 0]A_address0,
	output A_ce0,
	output A_we0,
	output [31 : 0]A_dout0,
	input [31 : 0]A_din0,
	output [11 : 0]A_address1,
	output A_ce1,
	output A_we1,
	output [31 : 0]A_dout1,
	input [31 : 0]A_din1,

	output [5 : 0]y1_address0,
	output y1_ce0,
	output y1_we0,
	output [31 : 0]y1_dout0,
	input [31 : 0]y1_din0,
	output [5 : 0]y1_address1,
	output y1_ce1,
	output y1_we1,
	output [31 : 0]y1_dout1,
	input [31 : 0]y1_din1,

	output [5 : 0]x2_address0,
	output x2_ce0,
	output x2_we0,
	output [31 : 0]x2_dout0,
	input [31 : 0]x2_din0,
	output [5 : 0]x2_address1,
	output x2_ce1,
	output x2_we1,
	output [31 : 0]x2_dout1,
	input [31 : 0]x2_din1,

	output [5 : 0]y2_address0,
	output y2_ce0,
	output y2_we0,
	output [31 : 0]y2_dout0,
	input [31 : 0]y2_din0,
	output [5 : 0]y2_address1,
	output y2_ce1,
	output y2_we1,
	output [31 : 0]y2_dout1,
	input [31 : 0]y2_din1

);

	wire phi_1_clk;
	wire phi_1_rst;
	wire [0 : 0]phi_1_in1_data;
	wire phi_1_in1_ready;
	wire phi_1_in1_valid;
	wire [5 : 0]phi_1_in2_data;
	wire phi_1_in2_ready;
	wire phi_1_in2_valid;
	wire [5 : 0]phi_1_in3_data;
	wire phi_1_in3_ready;
	wire phi_1_in3_valid;
	wire [5 : 0]phi_1_out1_data;
	wire phi_1_out1_ready;
	wire phi_1_out1_valid;

	wire load_4_clk;
	wire load_4_rst;
	wire [31 : 0]load_4_in1_data;
	wire load_4_in1_ready;
	wire load_4_in1_valid;
	wire [5 : 0]load_4_in2_data;
	wire load_4_in2_ready;
	wire load_4_in2_valid;
	wire [31 : 0]load_4_out1_data;
	wire load_4_out1_ready;
	wire load_4_out1_valid;
	wire [5 : 0]load_4_out2_data;
	wire load_4_out2_ready;
	wire load_4_out2_valid;

	wire brCst_block2_clk;
	wire brCst_block2_rst;
	wire [0 : 0]brCst_block2_in1_data;
	wire brCst_block2_in1_ready;
	wire brCst_block2_in1_valid;
	wire [0 : 0]brCst_block2_out1_data;
	wire brCst_block2_out1_ready;
	wire brCst_block2_out1_valid;

	wire cst_1_clk;
	wire cst_1_rst;
	wire [0 : 0]cst_1_in1_data;
	wire cst_1_in1_ready;
	wire cst_1_in1_valid;
	wire [0 : 0]cst_1_out1_data;
	wire cst_1_out1_ready;
	wire cst_1_out1_valid;

	wire fork_0_clk;
	wire fork_0_rst;
	wire [5 : 0]fork_0_in1_data;
	wire fork_0_in1_ready;
	wire fork_0_in1_valid;
	wire [5 : 0]fork_0_out1_data;
	wire fork_0_out1_ready;
	wire fork_0_out1_valid;
	wire [5 : 0]fork_0_out2_data;
	wire fork_0_out2_ready;
	wire fork_0_out2_valid;

	wire branch_1_clk;
	wire branch_1_rst;
	wire [31 : 0]branch_1_in1_data;
	wire branch_1_in1_ready;
	wire branch_1_in1_valid;
	wire [0 : 0]branch_1_in2_data;
	wire branch_1_in2_ready;
	wire branch_1_in2_valid;
	wire [31 : 0]branch_1_out1_data;
	wire branch_1_out1_ready;
	wire branch_1_out1_valid;
	wire [31 : 0]branch_1_out2_data;
	wire branch_1_out2_ready;
	wire branch_1_out2_valid;

	wire branch_2_clk;
	wire branch_2_rst;
	wire [0 : 0]branch_2_in1_data;
	wire branch_2_in1_ready;
	wire branch_2_in1_valid;
	wire [0 : 0]branch_2_in2_data;
	wire branch_2_in2_ready;
	wire branch_2_in2_valid;
	wire [0 : 0]branch_2_out1_data;
	wire branch_2_out1_ready;
	wire branch_2_out1_valid;
	wire [0 : 0]branch_2_out2_data;
	wire branch_2_out2_ready;
	wire branch_2_out2_valid;

	wire branch_3_clk;
	wire branch_3_rst;
	wire [5 : 0]branch_3_in1_data;
	wire branch_3_in1_ready;
	wire branch_3_in1_valid;
	wire [0 : 0]branch_3_in2_data;
	wire branch_3_in2_ready;
	wire branch_3_in2_valid;
	wire [5 : 0]branch_3_out1_data;
	wire branch_3_out1_ready;
	wire branch_3_out1_valid;
	wire [5 : 0]branch_3_out2_data;
	wire branch_3_out2_ready;
	wire branch_3_out2_valid;

	wire fork_15_clk;
	wire fork_15_rst;
	wire [0 : 0]fork_15_in1_data;
	wire fork_15_in1_ready;
	wire fork_15_in1_valid;
	wire [0 : 0]fork_15_out1_data;
	wire fork_15_out1_ready;
	wire fork_15_out1_valid;
	wire [0 : 0]fork_15_out2_data;
	wire fork_15_out2_ready;
	wire fork_15_out2_valid;
	wire [0 : 0]fork_15_out3_data;
	wire fork_15_out3_ready;
	wire fork_15_out3_valid;
	wire [0 : 0]fork_15_out4_data;
	wire fork_15_out4_ready;
	wire fork_15_out4_valid;

	wire phiC_6_clk;
	wire phiC_6_rst;
	wire [0 : 0]phiC_6_in1_data;
	wire phiC_6_in1_ready;
	wire phiC_6_in1_valid;
	wire [0 : 0]phiC_6_in2_data;
	wire phiC_6_in2_ready;
	wire phiC_6_in2_valid;
	wire [0 : 0]phiC_6_out1_data;
	wire phiC_6_out1_ready;
	wire phiC_6_out1_valid;
	wire [0 : 0]phiC_6_out2_data;
	wire phiC_6_out2_ready;
	wire phiC_6_out2_valid;

	wire forkC_25_clk;
	wire forkC_25_rst;
	wire [0 : 0]forkC_25_in1_data;
	wire forkC_25_in1_ready;
	wire forkC_25_in1_valid;
	wire [0 : 0]forkC_25_out1_data;
	wire forkC_25_out1_ready;
	wire forkC_25_out1_valid;
	wire [0 : 0]forkC_25_out2_data;
	wire forkC_25_out2_ready;
	wire forkC_25_out2_valid;
	wire [0 : 0]forkC_25_out3_data;
	wire forkC_25_out3_ready;
	wire forkC_25_out3_valid;

	wire branchC_17_clk;
	wire branchC_17_rst;
	wire [0 : 0]branchC_17_in1_data;
	wire branchC_17_in1_ready;
	wire branchC_17_in1_valid;
	wire [0 : 0]branchC_17_in2_data;
	wire branchC_17_in2_ready;
	wire branchC_17_in2_valid;
	wire [0 : 0]branchC_17_out1_data;
	wire branchC_17_out1_ready;
	wire branchC_17_out1_valid;
	wire [0 : 0]branchC_17_out2_data;
	wire branchC_17_out2_ready;
	wire branchC_17_out2_valid;

	wire brCst_block1_clk;
	wire brCst_block1_rst;
	wire [0 : 0]brCst_block1_in1_data;
	wire brCst_block1_in1_ready;
	wire brCst_block1_in1_valid;
	wire [0 : 0]brCst_block1_out1_data;
	wire brCst_block1_out1_ready;
	wire brCst_block1_out1_valid;

	wire cst_0_clk;
	wire cst_0_rst;
	wire [0 : 0]cst_0_in1_data;
	wire cst_0_in1_ready;
	wire cst_0_in1_valid;
	wire [0 : 0]cst_0_out1_data;
	wire cst_0_out1_ready;
	wire cst_0_out1_valid;

	wire branch_0_clk;
	wire branch_0_rst;
	wire [0 : 0]branch_0_in1_data;
	wire branch_0_in1_ready;
	wire branch_0_in1_valid;
	wire [0 : 0]branch_0_in2_data;
	wire branch_0_in2_ready;
	wire branch_0_in2_valid;
	wire [0 : 0]branch_0_out1_data;
	wire branch_0_out1_ready;
	wire branch_0_out1_valid;
	wire [0 : 0]branch_0_out2_data;
	wire branch_0_out2_ready;
	wire branch_0_out2_valid;

	wire start_0_clk;
	wire start_0_rst;
	wire [0 : 0]start_0_in1_data;
	wire start_0_in1_ready;
	wire start_0_in1_valid;
	wire [0 : 0]start_0_out1_data;
	wire start_0_out1_ready;
	wire start_0_out1_valid;

	wire forkC_23_clk;
	wire forkC_23_rst;
	wire [0 : 0]forkC_23_in1_data;
	wire forkC_23_in1_ready;
	wire forkC_23_in1_valid;
	wire [0 : 0]forkC_23_out1_data;
	wire forkC_23_out1_ready;
	wire forkC_23_out1_valid;
	wire [0 : 0]forkC_23_out2_data;
	wire forkC_23_out2_ready;
	wire forkC_23_out2_valid;
	wire [0 : 0]forkC_23_out3_data;
	wire forkC_23_out3_ready;
	wire forkC_23_out3_valid;

	wire branchC_16_clk;
	wire branchC_16_rst;
	wire [0 : 0]branchC_16_in1_data;
	wire branchC_16_in1_ready;
	wire branchC_16_in1_valid;
	wire [0 : 0]branchC_16_in2_data;
	wire branchC_16_in2_ready;
	wire branchC_16_in2_valid;
	wire [0 : 0]branchC_16_out1_data;
	wire branchC_16_out1_ready;
	wire branchC_16_out1_valid;
	wire [0 : 0]branchC_16_out2_data;
	wire branchC_16_out2_ready;
	wire branchC_16_out2_valid;

	wire fork_24_clk;
	wire fork_24_rst;
	wire [0 : 0]fork_24_in1_data;
	wire fork_24_in1_ready;
	wire fork_24_in1_valid;
	wire [0 : 0]fork_24_out1_data;
	wire fork_24_out1_ready;
	wire fork_24_out1_valid;
	wire [0 : 0]fork_24_out2_data;
	wire fork_24_out2_ready;
	wire fork_24_out2_valid;

	wire phi_27_clk;
	wire phi_27_rst;
	wire [0 : 0]phi_27_in1_data;
	wire phi_27_in1_ready;
	wire phi_27_in1_valid;
	wire [5 : 0]phi_27_in2_data;
	wire phi_27_in2_ready;
	wire phi_27_in2_valid;
	wire [5 : 0]phi_27_in3_data;
	wire phi_27_in3_ready;
	wire phi_27_in3_valid;
	wire [5 : 0]phi_27_out1_data;
	wire phi_27_out1_ready;
	wire phi_27_out1_valid;

	wire load_30_clk;
	wire load_30_rst;
	wire [31 : 0]load_30_in1_data;
	wire load_30_in1_ready;
	wire load_30_in1_valid;
	wire [5 : 0]load_30_in2_data;
	wire load_30_in2_ready;
	wire load_30_in2_valid;
	wire [31 : 0]load_30_out1_data;
	wire load_30_out1_ready;
	wire load_30_out1_valid;
	wire [5 : 0]load_30_out2_data;
	wire load_30_out2_ready;
	wire load_30_out2_valid;

	wire brCst_block6_clk;
	wire brCst_block6_rst;
	wire [0 : 0]brCst_block6_in1_data;
	wire brCst_block6_in1_ready;
	wire brCst_block6_in1_valid;
	wire [0 : 0]brCst_block6_out1_data;
	wire brCst_block6_out1_ready;
	wire brCst_block6_out1_valid;

	wire cst_8_clk;
	wire cst_8_rst;
	wire [0 : 0]cst_8_in1_data;
	wire cst_8_in1_ready;
	wire cst_8_in1_valid;
	wire [0 : 0]cst_8_out1_data;
	wire cst_8_out1_ready;
	wire cst_8_out1_valid;

	wire fork_5_clk;
	wire fork_5_rst;
	wire [5 : 0]fork_5_in1_data;
	wire fork_5_in1_ready;
	wire fork_5_in1_valid;
	wire [5 : 0]fork_5_out1_data;
	wire fork_5_out1_ready;
	wire fork_5_out1_valid;
	wire [5 : 0]fork_5_out2_data;
	wire fork_5_out2_ready;
	wire fork_5_out2_valid;

	wire branch_9_clk;
	wire branch_9_rst;
	wire [31 : 0]branch_9_in1_data;
	wire branch_9_in1_ready;
	wire branch_9_in1_valid;
	wire [0 : 0]branch_9_in2_data;
	wire branch_9_in2_ready;
	wire branch_9_in2_valid;
	wire [31 : 0]branch_9_out1_data;
	wire branch_9_out1_ready;
	wire branch_9_out1_valid;
	wire [31 : 0]branch_9_out2_data;
	wire branch_9_out2_ready;
	wire branch_9_out2_valid;

	wire branch_10_clk;
	wire branch_10_rst;
	wire [0 : 0]branch_10_in1_data;
	wire branch_10_in1_ready;
	wire branch_10_in1_valid;
	wire [0 : 0]branch_10_in2_data;
	wire branch_10_in2_ready;
	wire branch_10_in2_valid;
	wire [0 : 0]branch_10_out1_data;
	wire branch_10_out1_ready;
	wire branch_10_out1_valid;
	wire [0 : 0]branch_10_out2_data;
	wire branch_10_out2_ready;
	wire branch_10_out2_valid;

	wire branch_11_clk;
	wire branch_11_rst;
	wire [5 : 0]branch_11_in1_data;
	wire branch_11_in1_ready;
	wire branch_11_in1_valid;
	wire [0 : 0]branch_11_in2_data;
	wire branch_11_in2_ready;
	wire branch_11_in2_valid;
	wire [5 : 0]branch_11_out1_data;
	wire branch_11_out1_ready;
	wire branch_11_out1_valid;
	wire [5 : 0]branch_11_out2_data;
	wire branch_11_out2_ready;
	wire branch_11_out2_valid;

	wire fork_19_clk;
	wire fork_19_rst;
	wire [0 : 0]fork_19_in1_data;
	wire fork_19_in1_ready;
	wire fork_19_in1_valid;
	wire [0 : 0]fork_19_out1_data;
	wire fork_19_out1_ready;
	wire fork_19_out1_valid;
	wire [0 : 0]fork_19_out2_data;
	wire fork_19_out2_ready;
	wire fork_19_out2_valid;
	wire [0 : 0]fork_19_out3_data;
	wire fork_19_out3_ready;
	wire fork_19_out3_valid;
	wire [0 : 0]fork_19_out4_data;
	wire fork_19_out4_ready;
	wire fork_19_out4_valid;

	wire phiC_10_clk;
	wire phiC_10_rst;
	wire [0 : 0]phiC_10_in1_data;
	wire phiC_10_in1_ready;
	wire phiC_10_in1_valid;
	wire [0 : 0]phiC_10_in2_data;
	wire phiC_10_in2_ready;
	wire phiC_10_in2_valid;
	wire [0 : 0]phiC_10_out1_data;
	wire phiC_10_out1_ready;
	wire phiC_10_out1_valid;
	wire [0 : 0]phiC_10_out2_data;
	wire phiC_10_out2_ready;
	wire phiC_10_out2_valid;

	wire forkC_31_clk;
	wire forkC_31_rst;
	wire [0 : 0]forkC_31_in1_data;
	wire forkC_31_in1_ready;
	wire forkC_31_in1_valid;
	wire [0 : 0]forkC_31_out1_data;
	wire forkC_31_out1_ready;
	wire forkC_31_out1_valid;
	wire [0 : 0]forkC_31_out2_data;
	wire forkC_31_out2_ready;
	wire forkC_31_out2_valid;
	wire [0 : 0]forkC_31_out3_data;
	wire forkC_31_out3_ready;
	wire forkC_31_out3_valid;

	wire branchC_21_clk;
	wire branchC_21_rst;
	wire [0 : 0]branchC_21_in1_data;
	wire branchC_21_in1_ready;
	wire branchC_21_in1_valid;
	wire [0 : 0]branchC_21_in2_data;
	wire branchC_21_in2_ready;
	wire branchC_21_in2_valid;
	wire [0 : 0]branchC_21_out1_data;
	wire branchC_21_out1_ready;
	wire branchC_21_out1_valid;
	wire [0 : 0]branchC_21_out2_data;
	wire branchC_21_out2_ready;
	wire branchC_21_out2_valid;

	wire phi_32_clk;
	wire phi_32_rst;
	wire [0 : 0]phi_32_in1_data;
	wire phi_32_in1_ready;
	wire phi_32_in1_valid;
	wire [31 : 0]phi_32_in2_data;
	wire phi_32_in2_ready;
	wire phi_32_in2_valid;
	wire [31 : 0]phi_32_in3_data;
	wire phi_32_in3_ready;
	wire phi_32_in3_valid;
	wire [31 : 0]phi_32_out1_data;
	wire phi_32_out1_ready;
	wire phi_32_out1_valid;

	wire phi_33_clk;
	wire phi_33_rst;
	wire [0 : 0]phi_33_in1_data;
	wire phi_33_in1_ready;
	wire phi_33_in1_valid;
	wire [5 : 0]phi_33_in2_data;
	wire phi_33_in2_ready;
	wire phi_33_in2_valid;
	wire [5 : 0]phi_33_in3_data;
	wire phi_33_in3_ready;
	wire phi_33_in3_valid;
	wire [5 : 0]phi_33_out1_data;
	wire phi_33_out1_ready;
	wire phi_33_out1_valid;

	wire cst_9_clk;
	wire cst_9_rst;
	wire [2 : 0]cst_9_in1_data;
	wire cst_9_in1_ready;
	wire cst_9_in1_valid;
	wire [2 : 0]cst_9_out1_data;
	wire cst_9_out1_ready;
	wire cst_9_out1_valid;

	wire shl_34_clk;
	wire shl_34_rst;
	wire [10 : 0]shl_34_in1_data;
	wire shl_34_in1_ready;
	wire shl_34_in1_valid;
	wire [10 : 0]shl_34_in2_data;
	wire shl_34_in2_ready;
	wire shl_34_in2_valid;
	wire [10 : 0]shl_34_out1_data;
	wire shl_34_out1_ready;
	wire shl_34_out1_valid;

	wire add_35_clk;
	wire add_35_rst;
	wire [11 : 0]add_35_in1_data;
	wire add_35_in1_ready;
	wire add_35_in1_valid;
	wire [11 : 0]add_35_in2_data;
	wire add_35_in2_ready;
	wire add_35_in2_valid;
	wire [11 : 0]add_35_out1_data;
	wire add_35_out1_ready;
	wire add_35_out1_valid;

	wire load_38_clk;
	wire load_38_rst;
	wire [31 : 0]load_38_in1_data;
	wire load_38_in1_ready;
	wire load_38_in1_valid;
	wire [11 : 0]load_38_in2_data;
	wire load_38_in2_ready;
	wire load_38_in2_valid;
	wire [31 : 0]load_38_out1_data;
	wire load_38_out1_ready;
	wire load_38_out1_valid;
	wire [11 : 0]load_38_out2_data;
	wire load_38_out2_ready;
	wire load_38_out2_valid;

	wire load_41_clk;
	wire load_41_rst;
	wire [31 : 0]load_41_in1_data;
	wire load_41_in1_ready;
	wire load_41_in1_valid;
	wire [5 : 0]load_41_in2_data;
	wire load_41_in2_ready;
	wire load_41_in2_valid;
	wire [31 : 0]load_41_out1_data;
	wire load_41_out1_ready;
	wire load_41_out1_valid;
	wire [5 : 0]load_41_out2_data;
	wire load_41_out2_ready;
	wire load_41_out2_valid;

	wire cst_10_clk;
	wire cst_10_rst;
	wire [0 : 0]cst_10_in1_data;
	wire cst_10_in1_ready;
	wire cst_10_in1_valid;
	wire [0 : 0]cst_10_out1_data;
	wire cst_10_out1_ready;
	wire cst_10_out1_valid;

	wire add_44_clk;
	wire add_44_rst;
	wire [5 : 0]add_44_in1_data;
	wire add_44_in1_ready;
	wire add_44_in1_valid;
	wire [5 : 0]add_44_in2_data;
	wire add_44_in2_ready;
	wire add_44_in2_valid;
	wire [5 : 0]add_44_out1_data;
	wire add_44_out1_ready;
	wire add_44_out1_valid;

	wire cst_11_clk;
	wire cst_11_rst;
	wire [5 : 0]cst_11_in1_data;
	wire cst_11_in1_ready;
	wire cst_11_in1_valid;
	wire [5 : 0]cst_11_out1_data;
	wire cst_11_out1_ready;
	wire cst_11_out1_valid;

	wire icmp_45_clk;
	wire icmp_45_rst;
	wire [5 : 0]icmp_45_in1_data;
	wire icmp_45_in1_ready;
	wire icmp_45_in1_valid;
	wire [5 : 0]icmp_45_in2_data;
	wire icmp_45_in2_ready;
	wire icmp_45_in2_valid;
	wire [0 : 0]icmp_45_out1_data;
	wire icmp_45_out1_ready;
	wire icmp_45_out1_valid;

	wire phi_n5_clk;
	wire phi_n5_rst;
	wire [5 : 0]phi_n5_in1_data;
	wire phi_n5_in1_ready;
	wire phi_n5_in1_valid;
	wire [5 : 0]phi_n5_in2_data;
	wire phi_n5_in2_ready;
	wire phi_n5_in2_valid;
	wire [5 : 0]phi_n5_out1_data;
	wire phi_n5_out1_ready;
	wire phi_n5_out1_valid;

	wire fork_6_clk;
	wire fork_6_rst;
	wire [5 : 0]fork_6_in1_data;
	wire fork_6_in1_ready;
	wire fork_6_in1_valid;
	wire [5 : 0]fork_6_out1_data;
	wire fork_6_out1_ready;
	wire fork_6_out1_valid;
	wire [5 : 0]fork_6_out2_data;
	wire fork_6_out2_ready;
	wire fork_6_out2_valid;
	wire [5 : 0]fork_6_out3_data;
	wire fork_6_out3_ready;
	wire fork_6_out3_valid;

	wire fork_8_clk;
	wire fork_8_rst;
	wire [5 : 0]fork_8_in1_data;
	wire fork_8_in1_ready;
	wire fork_8_in1_valid;
	wire [5 : 0]fork_8_out1_data;
	wire fork_8_out1_ready;
	wire fork_8_out1_valid;
	wire [5 : 0]fork_8_out2_data;
	wire fork_8_out2_ready;
	wire fork_8_out2_valid;

	wire fork_13_clk;
	wire fork_13_rst;
	wire [5 : 0]fork_13_in1_data;
	wire fork_13_in1_ready;
	wire fork_13_in1_valid;
	wire [5 : 0]fork_13_out1_data;
	wire fork_13_out1_ready;
	wire fork_13_out1_valid;
	wire [5 : 0]fork_13_out2_data;
	wire fork_13_out2_ready;
	wire fork_13_out2_valid;

	wire branch_12_clk;
	wire branch_12_rst;
	wire [31 : 0]branch_12_in1_data;
	wire branch_12_in1_ready;
	wire branch_12_in1_valid;
	wire [0 : 0]branch_12_in2_data;
	wire branch_12_in2_ready;
	wire branch_12_in2_valid;
	wire [31 : 0]branch_12_out1_data;
	wire branch_12_out1_ready;
	wire branch_12_out1_valid;
	wire [31 : 0]branch_12_out2_data;
	wire branch_12_out2_ready;
	wire branch_12_out2_valid;

	wire branch_13_clk;
	wire branch_13_rst;
	wire [5 : 0]branch_13_in1_data;
	wire branch_13_in1_ready;
	wire branch_13_in1_valid;
	wire [0 : 0]branch_13_in2_data;
	wire branch_13_in2_ready;
	wire branch_13_in2_valid;
	wire [5 : 0]branch_13_out1_data;
	wire branch_13_out1_ready;
	wire branch_13_out1_valid;
	wire [5 : 0]branch_13_out2_data;
	wire branch_13_out2_ready;
	wire branch_13_out2_valid;

	wire branch_14_clk;
	wire branch_14_rst;
	wire [5 : 0]branch_14_in1_data;
	wire branch_14_in1_ready;
	wire branch_14_in1_valid;
	wire [0 : 0]branch_14_in2_data;
	wire branch_14_in2_ready;
	wire branch_14_in2_valid;
	wire [5 : 0]branch_14_out1_data;
	wire branch_14_out1_ready;
	wire branch_14_out1_valid;
	wire [5 : 0]branch_14_out2_data;
	wire branch_14_out2_ready;
	wire branch_14_out2_valid;

	wire fork_20_clk;
	wire fork_20_rst;
	wire [0 : 0]fork_20_in1_data;
	wire fork_20_in1_ready;
	wire fork_20_in1_valid;
	wire [0 : 0]fork_20_out1_data;
	wire fork_20_out1_ready;
	wire fork_20_out1_valid;
	wire [0 : 0]fork_20_out2_data;
	wire fork_20_out2_ready;
	wire fork_20_out2_valid;
	wire [0 : 0]fork_20_out3_data;
	wire fork_20_out3_ready;
	wire fork_20_out3_valid;
	wire [0 : 0]fork_20_out4_data;
	wire fork_20_out4_ready;
	wire fork_20_out4_valid;

	wire phiC_11_clk;
	wire phiC_11_rst;
	wire [0 : 0]phiC_11_in1_data;
	wire phiC_11_in1_ready;
	wire phiC_11_in1_valid;
	wire [0 : 0]phiC_11_in2_data;
	wire phiC_11_in2_ready;
	wire phiC_11_in2_valid;
	wire [0 : 0]phiC_11_out1_data;
	wire phiC_11_out1_ready;
	wire phiC_11_out1_valid;
	wire [0 : 0]phiC_11_out2_data;
	wire phiC_11_out2_ready;
	wire phiC_11_out2_valid;

	wire branchC_22_clk;
	wire branchC_22_rst;
	wire [0 : 0]branchC_22_in1_data;
	wire branchC_22_in1_ready;
	wire branchC_22_in1_valid;
	wire [0 : 0]branchC_22_in2_data;
	wire branchC_22_in2_ready;
	wire branchC_22_in2_valid;
	wire [0 : 0]branchC_22_out1_data;
	wire branchC_22_out1_ready;
	wire branchC_22_out1_valid;
	wire [0 : 0]branchC_22_out2_data;
	wire branchC_22_out2_ready;
	wire branchC_22_out2_valid;

	wire source_5_clk;
	wire source_5_rst;
	wire [2 : 0]source_5_out1_data;
	wire source_5_out1_ready;
	wire source_5_out1_valid;

	wire source_6_clk;
	wire source_6_rst;
	wire [0 : 0]source_6_out1_data;
	wire source_6_out1_ready;
	wire source_6_out1_valid;

	wire source_7_clk;
	wire source_7_rst;
	wire [5 : 0]source_7_out1_data;
	wire source_7_out1_ready;
	wire source_7_out1_valid;

	wire fork_39_clk;
	wire fork_39_rst;
	wire [0 : 0]fork_39_in1_data;
	wire fork_39_in1_ready;
	wire fork_39_in1_valid;
	wire [0 : 0]fork_39_out1_data;
	wire fork_39_out1_ready;
	wire fork_39_out1_valid;
	wire [0 : 0]fork_39_out2_data;
	wire fork_39_out2_ready;
	wire fork_39_out2_valid;

	wire store_1_clk;
	wire store_1_rst;
	wire [31 : 0]store_1_in1_data;
	wire store_1_in1_ready;
	wire store_1_in1_valid;
	wire [5 : 0]store_1_in2_data;
	wire store_1_in2_ready;
	wire store_1_in2_valid;
	wire [31 : 0]store_1_out1_data;
	wire store_1_out1_ready;
	wire store_1_out1_valid;
	wire [5 : 0]store_1_out2_data;
	wire store_1_out2_ready;
	wire store_1_out2_valid;

	wire cst_12_clk;
	wire cst_12_rst;
	wire [0 : 0]cst_12_in1_data;
	wire cst_12_in1_ready;
	wire cst_12_in1_valid;
	wire [0 : 0]cst_12_out1_data;
	wire cst_12_out1_ready;
	wire cst_12_out1_valid;

	wire add_49_clk;
	wire add_49_rst;
	wire [5 : 0]add_49_in1_data;
	wire add_49_in1_ready;
	wire add_49_in1_valid;
	wire [5 : 0]add_49_in2_data;
	wire add_49_in2_ready;
	wire add_49_in2_valid;
	wire [5 : 0]add_49_out1_data;
	wire add_49_out1_ready;
	wire add_49_out1_valid;

	wire cst_13_clk;
	wire cst_13_rst;
	wire [5 : 0]cst_13_in1_data;
	wire cst_13_in1_ready;
	wire cst_13_in1_valid;
	wire [5 : 0]cst_13_out1_data;
	wire cst_13_out1_ready;
	wire cst_13_out1_valid;

	wire icmp_50_clk;
	wire icmp_50_rst;
	wire [5 : 0]icmp_50_in1_data;
	wire icmp_50_in1_ready;
	wire icmp_50_in1_valid;
	wire [5 : 0]icmp_50_in2_data;
	wire icmp_50_in2_ready;
	wire icmp_50_in2_valid;
	wire [0 : 0]icmp_50_out1_data;
	wire icmp_50_out1_ready;
	wire icmp_50_out1_valid;

	wire phi_n3_clk;
	wire phi_n3_rst;
	wire [31 : 0]phi_n3_in1_data;
	wire phi_n3_in1_ready;
	wire phi_n3_in1_valid;
	wire [31 : 0]phi_n3_out1_data;
	wire phi_n3_out1_ready;
	wire phi_n3_out1_valid;

	wire phi_n4_clk;
	wire phi_n4_rst;
	wire [5 : 0]phi_n4_in1_data;
	wire phi_n4_in1_ready;
	wire phi_n4_in1_valid;
	wire [5 : 0]phi_n4_out1_data;
	wire phi_n4_out1_ready;
	wire phi_n4_out1_valid;

	wire fork_9_clk;
	wire fork_9_rst;
	wire [5 : 0]fork_9_in1_data;
	wire fork_9_in1_ready;
	wire fork_9_in1_valid;
	wire [5 : 0]fork_9_out1_data;
	wire fork_9_out1_ready;
	wire fork_9_out1_valid;
	wire [5 : 0]fork_9_out2_data;
	wire fork_9_out2_ready;
	wire fork_9_out2_valid;

	wire fork_12_clk;
	wire fork_12_rst;
	wire [5 : 0]fork_12_in1_data;
	wire fork_12_in1_ready;
	wire fork_12_in1_valid;
	wire [5 : 0]fork_12_out1_data;
	wire fork_12_out1_ready;
	wire fork_12_out1_valid;
	wire [5 : 0]fork_12_out2_data;
	wire fork_12_out2_ready;
	wire fork_12_out2_valid;

	wire branch_15_clk;
	wire branch_15_rst;
	wire [5 : 0]branch_15_in1_data;
	wire branch_15_in1_ready;
	wire branch_15_in1_valid;
	wire [0 : 0]branch_15_in2_data;
	wire branch_15_in2_ready;
	wire branch_15_in2_valid;
	wire [5 : 0]branch_15_out1_data;
	wire branch_15_out1_ready;
	wire branch_15_out1_valid;
	wire [5 : 0]branch_15_out2_data;
	wire branch_15_out2_ready;
	wire branch_15_out2_valid;

	wire cst_15_clk;
	wire cst_15_rst;
	wire [0 : 0]cst_15_in1_data;
	wire cst_15_in1_ready;
	wire cst_15_in1_valid;
	wire [0 : 0]cst_15_out1_data;
	wire cst_15_out1_ready;
	wire cst_15_out1_valid;

	wire phiC_12_clk;
	wire phiC_12_rst;
	wire [0 : 0]phiC_12_in1_data;
	wire phiC_12_in1_ready;
	wire phiC_12_in1_valid;
	wire [0 : 0]phiC_12_out1_data;
	wire phiC_12_out1_ready;
	wire phiC_12_out1_valid;

	wire forkC_33_clk;
	wire forkC_33_rst;
	wire [0 : 0]forkC_33_in1_data;
	wire forkC_33_in1_ready;
	wire forkC_33_in1_valid;
	wire [0 : 0]forkC_33_out1_data;
	wire forkC_33_out1_ready;
	wire forkC_33_out1_valid;
	wire [0 : 0]forkC_33_out2_data;
	wire forkC_33_out2_ready;
	wire forkC_33_out2_valid;

	wire branchC_23_clk;
	wire branchC_23_rst;
	wire [0 : 0]branchC_23_in1_data;
	wire branchC_23_in1_ready;
	wire branchC_23_in1_valid;
	wire [0 : 0]branchC_23_in2_data;
	wire branchC_23_in2_ready;
	wire branchC_23_in2_valid;
	wire [0 : 0]branchC_23_out1_data;
	wire branchC_23_out1_ready;
	wire branchC_23_out1_valid;
	wire [0 : 0]branchC_23_out2_data;
	wire branchC_23_out2_ready;
	wire branchC_23_out2_valid;

	wire fork_34_clk;
	wire fork_34_rst;
	wire [0 : 0]fork_34_in1_data;
	wire fork_34_in1_ready;
	wire fork_34_in1_valid;
	wire [0 : 0]fork_34_out1_data;
	wire fork_34_out1_ready;
	wire fork_34_out1_valid;
	wire [0 : 0]fork_34_out2_data;
	wire fork_34_out2_ready;
	wire fork_34_out2_valid;

	wire source_8_clk;
	wire source_8_rst;
	wire [0 : 0]source_8_out1_data;
	wire source_8_out1_ready;
	wire source_8_out1_valid;

	wire source_9_clk;
	wire source_9_rst;
	wire [5 : 0]source_9_out1_data;
	wire source_9_out1_ready;
	wire source_9_out1_valid;

	wire brCst_block5_clk;
	wire brCst_block5_rst;
	wire [0 : 0]brCst_block5_in1_data;
	wire brCst_block5_in1_ready;
	wire brCst_block5_in1_valid;
	wire [0 : 0]brCst_block5_out1_data;
	wire brCst_block5_out1_ready;
	wire brCst_block5_out1_valid;

	wire cst_7_clk;
	wire cst_7_rst;
	wire [0 : 0]cst_7_in1_data;
	wire cst_7_in1_ready;
	wire cst_7_in1_valid;
	wire [0 : 0]cst_7_out1_data;
	wire cst_7_out1_ready;
	wire cst_7_out1_valid;

	wire branch_8_clk;
	wire branch_8_rst;
	wire [0 : 0]branch_8_in1_data;
	wire branch_8_in1_ready;
	wire branch_8_in1_valid;
	wire [0 : 0]branch_8_in2_data;
	wire branch_8_in2_ready;
	wire branch_8_in2_valid;
	wire [0 : 0]branch_8_out1_data;
	wire branch_8_out1_ready;
	wire branch_8_out1_valid;
	wire [0 : 0]branch_8_out2_data;
	wire branch_8_out2_ready;
	wire branch_8_out2_valid;

	wire phiC_9_clk;
	wire phiC_9_rst;
	wire [0 : 0]phiC_9_in1_data;
	wire phiC_9_in1_ready;
	wire phiC_9_in1_valid;
	wire [0 : 0]phiC_9_out1_data;
	wire phiC_9_out1_ready;
	wire phiC_9_out1_valid;

	wire forkC_29_clk;
	wire forkC_29_rst;
	wire [0 : 0]forkC_29_in1_data;
	wire forkC_29_in1_ready;
	wire forkC_29_in1_valid;
	wire [0 : 0]forkC_29_out1_data;
	wire forkC_29_out1_ready;
	wire forkC_29_out1_valid;
	wire [0 : 0]forkC_29_out2_data;
	wire forkC_29_out2_ready;
	wire forkC_29_out2_valid;
	wire [0 : 0]forkC_29_out3_data;
	wire forkC_29_out3_ready;
	wire forkC_29_out3_valid;

	wire branchC_20_clk;
	wire branchC_20_rst;
	wire [0 : 0]branchC_20_in1_data;
	wire branchC_20_in1_ready;
	wire branchC_20_in1_valid;
	wire [0 : 0]branchC_20_in2_data;
	wire branchC_20_in2_ready;
	wire branchC_20_in2_valid;
	wire [0 : 0]branchC_20_out1_data;
	wire branchC_20_out1_ready;
	wire branchC_20_out1_valid;
	wire [0 : 0]branchC_20_out2_data;
	wire branchC_20_out2_ready;
	wire branchC_20_out2_valid;

	wire fork_30_clk;
	wire fork_30_rst;
	wire [0 : 0]fork_30_in1_data;
	wire fork_30_in1_ready;
	wire fork_30_in1_valid;
	wire [0 : 0]fork_30_out1_data;
	wire fork_30_out1_ready;
	wire fork_30_out1_valid;
	wire [0 : 0]fork_30_out2_data;
	wire fork_30_out2_ready;
	wire fork_30_out2_valid;

	wire phi_6_clk;
	wire phi_6_rst;
	wire [0 : 0]phi_6_in1_data;
	wire phi_6_in1_ready;
	wire phi_6_in1_valid;
	wire [31 : 0]phi_6_in2_data;
	wire phi_6_in2_ready;
	wire phi_6_in2_valid;
	wire [31 : 0]phi_6_in3_data;
	wire phi_6_in3_ready;
	wire phi_6_in3_valid;
	wire [31 : 0]phi_6_out1_data;
	wire phi_6_out1_ready;
	wire phi_6_out1_valid;

	wire phi_7_clk;
	wire phi_7_rst;
	wire [0 : 0]phi_7_in1_data;
	wire phi_7_in1_ready;
	wire phi_7_in1_valid;
	wire [5 : 0]phi_7_in2_data;
	wire phi_7_in2_ready;
	wire phi_7_in2_valid;
	wire [5 : 0]phi_7_in3_data;
	wire phi_7_in3_ready;
	wire phi_7_in3_valid;
	wire [5 : 0]phi_7_out1_data;
	wire phi_7_out1_ready;
	wire phi_7_out1_valid;

	wire cst_2_clk;
	wire cst_2_rst;
	wire [2 : 0]cst_2_in1_data;
	wire cst_2_in1_ready;
	wire cst_2_in1_valid;
	wire [2 : 0]cst_2_out1_data;
	wire cst_2_out1_ready;
	wire cst_2_out1_valid;

	wire shl_8_clk;
	wire shl_8_rst;
	wire [10 : 0]shl_8_in1_data;
	wire shl_8_in1_ready;
	wire shl_8_in1_valid;
	wire [10 : 0]shl_8_in2_data;
	wire shl_8_in2_ready;
	wire shl_8_in2_valid;
	wire [10 : 0]shl_8_out1_data;
	wire shl_8_out1_ready;
	wire shl_8_out1_valid;

	wire add_9_clk;
	wire add_9_rst;
	wire [11 : 0]add_9_in1_data;
	wire add_9_in1_ready;
	wire add_9_in1_valid;
	wire [11 : 0]add_9_in2_data;
	wire add_9_in2_ready;
	wire add_9_in2_valid;
	wire [11 : 0]add_9_out1_data;
	wire add_9_out1_ready;
	wire add_9_out1_valid;

	wire load_12_clk;
	wire load_12_rst;
	wire [31 : 0]load_12_in1_data;
	wire load_12_in1_ready;
	wire load_12_in1_valid;
	wire [11 : 0]load_12_in2_data;
	wire load_12_in2_ready;
	wire load_12_in2_valid;
	wire [31 : 0]load_12_out1_data;
	wire load_12_out1_ready;
	wire load_12_out1_valid;
	wire [11 : 0]load_12_out2_data;
	wire load_12_out2_ready;
	wire load_12_out2_valid;

	wire load_15_clk;
	wire load_15_rst;
	wire [31 : 0]load_15_in1_data;
	wire load_15_in1_ready;
	wire load_15_in1_valid;
	wire [5 : 0]load_15_in2_data;
	wire load_15_in2_ready;
	wire load_15_in2_valid;
	wire [31 : 0]load_15_out1_data;
	wire load_15_out1_ready;
	wire load_15_out1_valid;
	wire [5 : 0]load_15_out2_data;
	wire load_15_out2_ready;
	wire load_15_out2_valid;

	wire cst_3_clk;
	wire cst_3_rst;
	wire [0 : 0]cst_3_in1_data;
	wire cst_3_in1_ready;
	wire cst_3_in1_valid;
	wire [0 : 0]cst_3_out1_data;
	wire cst_3_out1_ready;
	wire cst_3_out1_valid;

	wire add_18_clk;
	wire add_18_rst;
	wire [5 : 0]add_18_in1_data;
	wire add_18_in1_ready;
	wire add_18_in1_valid;
	wire [5 : 0]add_18_in2_data;
	wire add_18_in2_ready;
	wire add_18_in2_valid;
	wire [5 : 0]add_18_out1_data;
	wire add_18_out1_ready;
	wire add_18_out1_valid;

	wire cst_4_clk;
	wire cst_4_rst;
	wire [5 : 0]cst_4_in1_data;
	wire cst_4_in1_ready;
	wire cst_4_in1_valid;
	wire [5 : 0]cst_4_out1_data;
	wire cst_4_out1_ready;
	wire cst_4_out1_valid;

	wire icmp_19_clk;
	wire icmp_19_rst;
	wire [5 : 0]icmp_19_in1_data;
	wire icmp_19_in1_ready;
	wire icmp_19_in1_valid;
	wire [5 : 0]icmp_19_in2_data;
	wire icmp_19_in2_ready;
	wire icmp_19_in2_valid;
	wire [0 : 0]icmp_19_out1_data;
	wire icmp_19_out1_ready;
	wire icmp_19_out1_valid;

	wire phi_n2_clk;
	wire phi_n2_rst;
	wire [5 : 0]phi_n2_in1_data;
	wire phi_n2_in1_ready;
	wire phi_n2_in1_valid;
	wire [5 : 0]phi_n2_in2_data;
	wire phi_n2_in2_ready;
	wire phi_n2_in2_valid;
	wire [5 : 0]phi_n2_out1_data;
	wire phi_n2_out1_ready;
	wire phi_n2_out1_valid;

	wire fork_1_clk;
	wire fork_1_rst;
	wire [5 : 0]fork_1_in1_data;
	wire fork_1_in1_ready;
	wire fork_1_in1_valid;
	wire [5 : 0]fork_1_out1_data;
	wire fork_1_out1_ready;
	wire fork_1_out1_valid;
	wire [5 : 0]fork_1_out2_data;
	wire fork_1_out2_ready;
	wire fork_1_out2_valid;
	wire [5 : 0]fork_1_out3_data;
	wire fork_1_out3_ready;
	wire fork_1_out3_valid;

	wire fork_3_clk;
	wire fork_3_rst;
	wire [5 : 0]fork_3_in1_data;
	wire fork_3_in1_ready;
	wire fork_3_in1_valid;
	wire [5 : 0]fork_3_out1_data;
	wire fork_3_out1_ready;
	wire fork_3_out1_valid;
	wire [5 : 0]fork_3_out2_data;
	wire fork_3_out2_ready;
	wire fork_3_out2_valid;

	wire fork_11_clk;
	wire fork_11_rst;
	wire [5 : 0]fork_11_in1_data;
	wire fork_11_in1_ready;
	wire fork_11_in1_valid;
	wire [5 : 0]fork_11_out1_data;
	wire fork_11_out1_ready;
	wire fork_11_out1_valid;
	wire [5 : 0]fork_11_out2_data;
	wire fork_11_out2_ready;
	wire fork_11_out2_valid;

	wire branch_4_clk;
	wire branch_4_rst;
	wire [31 : 0]branch_4_in1_data;
	wire branch_4_in1_ready;
	wire branch_4_in1_valid;
	wire [0 : 0]branch_4_in2_data;
	wire branch_4_in2_ready;
	wire branch_4_in2_valid;
	wire [31 : 0]branch_4_out1_data;
	wire branch_4_out1_ready;
	wire branch_4_out1_valid;
	wire [31 : 0]branch_4_out2_data;
	wire branch_4_out2_ready;
	wire branch_4_out2_valid;

	wire branch_5_clk;
	wire branch_5_rst;
	wire [5 : 0]branch_5_in1_data;
	wire branch_5_in1_ready;
	wire branch_5_in1_valid;
	wire [0 : 0]branch_5_in2_data;
	wire branch_5_in2_ready;
	wire branch_5_in2_valid;
	wire [5 : 0]branch_5_out1_data;
	wire branch_5_out1_ready;
	wire branch_5_out1_valid;
	wire [5 : 0]branch_5_out2_data;
	wire branch_5_out2_ready;
	wire branch_5_out2_valid;

	wire branch_6_clk;
	wire branch_6_rst;
	wire [5 : 0]branch_6_in1_data;
	wire branch_6_in1_ready;
	wire branch_6_in1_valid;
	wire [0 : 0]branch_6_in2_data;
	wire branch_6_in2_ready;
	wire branch_6_in2_valid;
	wire [5 : 0]branch_6_out1_data;
	wire branch_6_out1_ready;
	wire branch_6_out1_valid;
	wire [5 : 0]branch_6_out2_data;
	wire branch_6_out2_ready;
	wire branch_6_out2_valid;

	wire fork_16_clk;
	wire fork_16_rst;
	wire [0 : 0]fork_16_in1_data;
	wire fork_16_in1_ready;
	wire fork_16_in1_valid;
	wire [0 : 0]fork_16_out1_data;
	wire fork_16_out1_ready;
	wire fork_16_out1_valid;
	wire [0 : 0]fork_16_out2_data;
	wire fork_16_out2_ready;
	wire fork_16_out2_valid;
	wire [0 : 0]fork_16_out3_data;
	wire fork_16_out3_ready;
	wire fork_16_out3_valid;
	wire [0 : 0]fork_16_out4_data;
	wire fork_16_out4_ready;
	wire fork_16_out4_valid;

	wire phiC_7_clk;
	wire phiC_7_rst;
	wire [0 : 0]phiC_7_in1_data;
	wire phiC_7_in1_ready;
	wire phiC_7_in1_valid;
	wire [0 : 0]phiC_7_in2_data;
	wire phiC_7_in2_ready;
	wire phiC_7_in2_valid;
	wire [0 : 0]phiC_7_out1_data;
	wire phiC_7_out1_ready;
	wire phiC_7_out1_valid;
	wire [0 : 0]phiC_7_out2_data;
	wire phiC_7_out2_ready;
	wire phiC_7_out2_valid;

	wire branchC_18_clk;
	wire branchC_18_rst;
	wire [0 : 0]branchC_18_in1_data;
	wire branchC_18_in1_ready;
	wire branchC_18_in1_valid;
	wire [0 : 0]branchC_18_in2_data;
	wire branchC_18_in2_ready;
	wire branchC_18_in2_valid;
	wire [0 : 0]branchC_18_out1_data;
	wire branchC_18_out1_ready;
	wire branchC_18_out1_valid;
	wire [0 : 0]branchC_18_out2_data;
	wire branchC_18_out2_ready;
	wire branchC_18_out2_valid;

	wire source_0_clk;
	wire source_0_rst;
	wire [2 : 0]source_0_out1_data;
	wire source_0_out1_ready;
	wire source_0_out1_valid;

	wire source_1_clk;
	wire source_1_rst;
	wire [0 : 0]source_1_out1_data;
	wire source_1_out1_ready;
	wire source_1_out1_valid;

	wire source_2_clk;
	wire source_2_rst;
	wire [5 : 0]source_2_out1_data;
	wire source_2_out1_ready;
	wire source_2_out1_valid;

	wire fork_37_clk;
	wire fork_37_rst;
	wire [0 : 0]fork_37_in1_data;
	wire fork_37_in1_ready;
	wire fork_37_in1_valid;
	wire [0 : 0]fork_37_out1_data;
	wire fork_37_out1_ready;
	wire fork_37_out1_valid;
	wire [0 : 0]fork_37_out2_data;
	wire fork_37_out2_ready;
	wire fork_37_out2_valid;

	wire store_0_clk;
	wire store_0_rst;
	wire [31 : 0]store_0_in1_data;
	wire store_0_in1_ready;
	wire store_0_in1_valid;
	wire [5 : 0]store_0_in2_data;
	wire store_0_in2_ready;
	wire store_0_in2_valid;
	wire [31 : 0]store_0_out1_data;
	wire store_0_out1_ready;
	wire store_0_out1_valid;
	wire [5 : 0]store_0_out2_data;
	wire store_0_out2_ready;
	wire store_0_out2_valid;

	wire cst_5_clk;
	wire cst_5_rst;
	wire [0 : 0]cst_5_in1_data;
	wire cst_5_in1_ready;
	wire cst_5_in1_valid;
	wire [0 : 0]cst_5_out1_data;
	wire cst_5_out1_ready;
	wire cst_5_out1_valid;

	wire add_23_clk;
	wire add_23_rst;
	wire [5 : 0]add_23_in1_data;
	wire add_23_in1_ready;
	wire add_23_in1_valid;
	wire [5 : 0]add_23_in2_data;
	wire add_23_in2_ready;
	wire add_23_in2_valid;
	wire [5 : 0]add_23_out1_data;
	wire add_23_out1_ready;
	wire add_23_out1_valid;

	wire cst_6_clk;
	wire cst_6_rst;
	wire [5 : 0]cst_6_in1_data;
	wire cst_6_in1_ready;
	wire cst_6_in1_valid;
	wire [5 : 0]cst_6_out1_data;
	wire cst_6_out1_ready;
	wire cst_6_out1_valid;

	wire icmp_24_clk;
	wire icmp_24_rst;
	wire [5 : 0]icmp_24_in1_data;
	wire icmp_24_in1_ready;
	wire icmp_24_in1_valid;
	wire [5 : 0]icmp_24_in2_data;
	wire icmp_24_in2_ready;
	wire icmp_24_in2_valid;
	wire [0 : 0]icmp_24_out1_data;
	wire icmp_24_out1_ready;
	wire icmp_24_out1_valid;

	wire phi_n0_clk;
	wire phi_n0_rst;
	wire [31 : 0]phi_n0_in1_data;
	wire phi_n0_in1_ready;
	wire phi_n0_in1_valid;
	wire [31 : 0]phi_n0_out1_data;
	wire phi_n0_out1_ready;
	wire phi_n0_out1_valid;

	wire phi_n1_clk;
	wire phi_n1_rst;
	wire [5 : 0]phi_n1_in1_data;
	wire phi_n1_in1_ready;
	wire phi_n1_in1_valid;
	wire [5 : 0]phi_n1_out1_data;
	wire phi_n1_out1_ready;
	wire phi_n1_out1_valid;

	wire fork_4_clk;
	wire fork_4_rst;
	wire [5 : 0]fork_4_in1_data;
	wire fork_4_in1_ready;
	wire fork_4_in1_valid;
	wire [5 : 0]fork_4_out1_data;
	wire fork_4_out1_ready;
	wire fork_4_out1_valid;
	wire [5 : 0]fork_4_out2_data;
	wire fork_4_out2_ready;
	wire fork_4_out2_valid;

	wire fork_10_clk;
	wire fork_10_rst;
	wire [5 : 0]fork_10_in1_data;
	wire fork_10_in1_ready;
	wire fork_10_in1_valid;
	wire [5 : 0]fork_10_out1_data;
	wire fork_10_out1_ready;
	wire fork_10_out1_valid;
	wire [5 : 0]fork_10_out2_data;
	wire fork_10_out2_ready;
	wire fork_10_out2_valid;

	wire branch_7_clk;
	wire branch_7_rst;
	wire [5 : 0]branch_7_in1_data;
	wire branch_7_in1_ready;
	wire branch_7_in1_valid;
	wire [0 : 0]branch_7_in2_data;
	wire branch_7_in2_ready;
	wire branch_7_in2_valid;
	wire [5 : 0]branch_7_out1_data;
	wire branch_7_out1_ready;
	wire branch_7_out1_valid;
	wire [5 : 0]branch_7_out2_data;
	wire branch_7_out2_ready;
	wire branch_7_out2_valid;

	wire cst_14_clk;
	wire cst_14_rst;
	wire [0 : 0]cst_14_in1_data;
	wire cst_14_in1_ready;
	wire cst_14_in1_valid;
	wire [0 : 0]cst_14_out1_data;
	wire cst_14_out1_ready;
	wire cst_14_out1_valid;

	wire phiC_8_clk;
	wire phiC_8_rst;
	wire [0 : 0]phiC_8_in1_data;
	wire phiC_8_in1_ready;
	wire phiC_8_in1_valid;
	wire [0 : 0]phiC_8_out1_data;
	wire phiC_8_out1_ready;
	wire phiC_8_out1_valid;

	wire forkC_27_clk;
	wire forkC_27_rst;
	wire [0 : 0]forkC_27_in1_data;
	wire forkC_27_in1_ready;
	wire forkC_27_in1_valid;
	wire [0 : 0]forkC_27_out1_data;
	wire forkC_27_out1_ready;
	wire forkC_27_out1_valid;
	wire [0 : 0]forkC_27_out2_data;
	wire forkC_27_out2_ready;
	wire forkC_27_out2_valid;

	wire branchC_19_clk;
	wire branchC_19_rst;
	wire [0 : 0]branchC_19_in1_data;
	wire branchC_19_in1_ready;
	wire branchC_19_in1_valid;
	wire [0 : 0]branchC_19_in2_data;
	wire branchC_19_in2_ready;
	wire branchC_19_in2_valid;
	wire [0 : 0]branchC_19_out1_data;
	wire branchC_19_out1_ready;
	wire branchC_19_out1_valid;
	wire [0 : 0]branchC_19_out2_data;
	wire branchC_19_out2_ready;
	wire branchC_19_out2_valid;

	wire fork_28_clk;
	wire fork_28_rst;
	wire [0 : 0]fork_28_in1_data;
	wire fork_28_in1_ready;
	wire fork_28_in1_valid;
	wire [0 : 0]fork_28_out1_data;
	wire fork_28_out1_ready;
	wire fork_28_out1_valid;
	wire [0 : 0]fork_28_out2_data;
	wire fork_28_out2_ready;
	wire fork_28_out2_valid;

	wire source_3_clk;
	wire source_3_rst;
	wire [0 : 0]source_3_out1_data;
	wire source_3_out1_ready;
	wire source_3_out1_valid;

	wire source_4_clk;
	wire source_4_rst;
	wire [5 : 0]source_4_out1_data;
	wire source_4_out1_ready;
	wire source_4_out1_valid;

	wire ret_0_clk;
	wire ret_0_rst;
	wire [0 : 0]ret_0_in1_data;
	wire ret_0_in1_ready;
	wire ret_0_in1_valid;
	wire [0 : 0]ret_0_out1_data;
	wire ret_0_out1_ready;
	wire ret_0_out1_valid;

	wire end_0_clk;
	wire end_0_rst;
	wire [0 : 0]end_0_in1_data;
	wire end_0_in1_ready;
	wire end_0_in1_valid;
	wire [0 : 0]end_0_in2_data;
	wire end_0_in2_ready;
	wire end_0_in2_valid;
	wire [0 : 0]end_0_in3_data;
	wire end_0_in3_ready;
	wire end_0_in3_valid;
	wire [0 : 0]end_0_in4_data;
	wire end_0_in4_ready;
	wire end_0_in4_valid;
	wire [0 : 0]end_0_in5_data;
	wire end_0_in5_ready;
	wire end_0_in5_valid;
	wire [0 : 0]end_0_in6_data;
	wire end_0_in6_ready;
	wire end_0_in6_valid;
	wire [0 : 0]end_0_out1_data;
	wire end_0_out1_ready;
	wire end_0_out1_valid;

	wire phiC_13_clk;
	wire phiC_13_rst;
	wire [0 : 0]phiC_13_in1_data;
	wire phiC_13_in1_ready;
	wire phiC_13_in1_valid;
	wire [0 : 0]phiC_13_out1_data;
	wire phiC_13_out1_ready;
	wire phiC_13_out1_valid;

	wire MC_x1_clk;
	wire MC_x1_rst;
	wire [31 : 0]MC_x1_in1_data;
	wire MC_x1_in1_ready;
	wire MC_x1_in1_valid;
	wire [5 : 0]MC_x1_in2_data;
	wire MC_x1_in2_ready;
	wire MC_x1_in2_valid;
	wire [5 : 0]MC_x1_in3_data;
	wire MC_x1_in3_ready;
	wire MC_x1_in3_valid;
	wire [31 : 0]MC_x1_in4_data;
	wire MC_x1_in4_ready;
	wire MC_x1_in4_valid;
	wire [31 : 0]MC_x1_out1_data;
	wire MC_x1_out1_ready;
	wire MC_x1_out1_valid;
	wire [0 : 0]MC_x1_out2_data;
	wire MC_x1_out2_ready;
	wire MC_x1_out2_valid;

	wire MC_A_clk;
	wire MC_A_rst;
	wire [11 : 0]MC_A_in1_data;
	wire MC_A_in1_ready;
	wire MC_A_in1_valid;
	wire [11 : 0]MC_A_in2_data;
	wire MC_A_in2_ready;
	wire MC_A_in2_valid;
	wire [31 : 0]MC_A_in3_data;
	wire MC_A_in3_ready;
	wire MC_A_in3_valid;
	wire [11 : 0]MC_A_in4_data;
	wire MC_A_in4_ready;
	wire MC_A_in4_valid;
	wire [31 : 0]MC_A_in5_data;
	wire MC_A_in5_ready;
	wire MC_A_in5_valid;
	wire [31 : 0]MC_A_out1_data;
	wire MC_A_out1_ready;
	wire MC_A_out1_valid;
	wire [31 : 0]MC_A_out2_data;
	wire MC_A_out2_ready;
	wire MC_A_out2_valid;
	wire [0 : 0]MC_A_out3_data;
	wire MC_A_out3_ready;
	wire MC_A_out3_valid;

	wire MC_y1_clk;
	wire MC_y1_rst;
	wire [5 : 0]MC_y1_in1_data;
	wire MC_y1_in1_ready;
	wire MC_y1_in1_valid;
	wire [31 : 0]MC_y1_in2_data;
	wire MC_y1_in2_ready;
	wire MC_y1_in2_valid;
	wire [5 : 0]MC_y1_in3_data;
	wire MC_y1_in3_ready;
	wire MC_y1_in3_valid;
	wire [31 : 0]MC_y1_in4_data;
	wire MC_y1_in4_ready;
	wire MC_y1_in4_valid;
	wire [31 : 0]MC_y1_out1_data;
	wire MC_y1_out1_ready;
	wire MC_y1_out1_valid;
	wire [0 : 0]MC_y1_out2_data;
	wire MC_y1_out2_ready;
	wire MC_y1_out2_valid;

	wire MC_x2_clk;
	wire MC_x2_rst;
	wire [31 : 0]MC_x2_in1_data;
	wire MC_x2_in1_ready;
	wire MC_x2_in1_valid;
	wire [5 : 0]MC_x2_in2_data;
	wire MC_x2_in2_ready;
	wire MC_x2_in2_valid;
	wire [5 : 0]MC_x2_in3_data;
	wire MC_x2_in3_ready;
	wire MC_x2_in3_valid;
	wire [31 : 0]MC_x2_in4_data;
	wire MC_x2_in4_ready;
	wire MC_x2_in4_valid;
	wire [31 : 0]MC_x2_out1_data;
	wire MC_x2_out1_ready;
	wire MC_x2_out1_valid;
	wire [0 : 0]MC_x2_out2_data;
	wire MC_x2_out2_ready;
	wire MC_x2_out2_valid;

	wire MC_y2_clk;
	wire MC_y2_rst;
	wire [5 : 0]MC_y2_in1_data;
	wire MC_y2_in1_ready;
	wire MC_y2_in1_valid;
	wire [31 : 0]MC_y2_in2_data;
	wire MC_y2_in2_ready;
	wire MC_y2_in2_valid;
	wire [5 : 0]MC_y2_in3_data;
	wire MC_y2_in3_ready;
	wire MC_y2_in3_valid;
	wire [31 : 0]MC_y2_in4_data;
	wire MC_y2_in4_ready;
	wire MC_y2_in4_valid;
	wire [31 : 0]MC_y2_out1_data;
	wire MC_y2_out1_ready;
	wire MC_y2_out1_valid;
	wire [0 : 0]MC_y2_out2_data;
	wire MC_y2_out2_ready;
	wire MC_y2_out2_valid;

	wire sink_0_clk;
	wire sink_0_rst;
	wire [0 : 0]sink_0_in1_data;
	wire sink_0_in1_ready;
	wire sink_0_in1_valid;

	wire sink_1_clk;
	wire sink_1_rst;
	wire [31 : 0]sink_1_in1_data;
	wire sink_1_in1_ready;
	wire sink_1_in1_valid;

	wire sink_2_clk;
	wire sink_2_rst;
	wire [0 : 0]sink_2_in1_data;
	wire sink_2_in1_ready;
	wire sink_2_in1_valid;

	wire sink_3_clk;
	wire sink_3_rst;
	wire [5 : 0]sink_3_in1_data;
	wire sink_3_in1_ready;
	wire sink_3_in1_valid;

	wire sink_4_clk;
	wire sink_4_rst;
	wire [5 : 0]sink_4_in1_data;
	wire sink_4_in1_ready;
	wire sink_4_in1_valid;

	wire sink_5_clk;
	wire sink_5_rst;
	wire [5 : 0]sink_5_in1_data;
	wire sink_5_in1_ready;
	wire sink_5_in1_valid;

	wire sink_6_clk;
	wire sink_6_rst;
	wire [0 : 0]sink_6_in1_data;
	wire sink_6_in1_ready;
	wire sink_6_in1_valid;

	wire sink_7_clk;
	wire sink_7_rst;
	wire [31 : 0]sink_7_in1_data;
	wire sink_7_in1_ready;
	wire sink_7_in1_valid;

	wire sink_8_clk;
	wire sink_8_rst;
	wire [0 : 0]sink_8_in1_data;
	wire sink_8_in1_ready;
	wire sink_8_in1_valid;

	wire sink_9_clk;
	wire sink_9_rst;
	wire [5 : 0]sink_9_in1_data;
	wire sink_9_in1_ready;
	wire sink_9_in1_valid;

	wire sink_10_clk;
	wire sink_10_rst;
	wire [5 : 0]sink_10_in1_data;
	wire sink_10_in1_ready;
	wire sink_10_in1_valid;

	wire sink_11_clk;
	wire sink_11_rst;
	wire [5 : 0]sink_11_in1_data;
	wire sink_11_in1_ready;
	wire sink_11_in1_valid;

	wire sink_12_clk;
	wire sink_12_rst;
	wire [0 : 0]sink_12_in1_data;
	wire sink_12_in1_ready;
	wire sink_12_in1_valid;

	wire sink_13_clk;
	wire sink_13_rst;
	wire [0 : 0]sink_13_in1_data;
	wire sink_13_in1_ready;
	wire sink_13_in1_valid;

	wire sink_14_clk;
	wire sink_14_rst;
	wire [0 : 0]sink_14_in1_data;
	wire sink_14_in1_ready;
	wire sink_14_in1_valid;

	wire sink_15_clk;
	wire sink_15_rst;
	wire [0 : 0]sink_15_in1_data;
	wire sink_15_in1_ready;
	wire sink_15_in1_valid;

	wire Buffer_100_clk;
	wire Buffer_100_rst;
	wire [31 : 0]Buffer_100_in1_data;
	wire Buffer_100_in1_ready;
	wire Buffer_100_in1_valid;
	wire [31 : 0]Buffer_100_out1_data;
	wire Buffer_100_out1_ready;
	wire Buffer_100_out1_valid;

	wire Buffer_101_clk;
	wire Buffer_101_rst;
	wire [31 : 0]Buffer_101_in1_data;
	wire Buffer_101_in1_ready;
	wire Buffer_101_in1_valid;
	wire [31 : 0]Buffer_101_out1_data;
	wire Buffer_101_out1_ready;
	wire Buffer_101_out1_valid;

	wire Buffer_102_clk;
	wire Buffer_102_rst;
	wire [31 : 0]Buffer_102_in1_data;
	wire Buffer_102_in1_ready;
	wire Buffer_102_in1_valid;
	wire [31 : 0]Buffer_102_out1_data;
	wire Buffer_102_out1_ready;
	wire Buffer_102_out1_valid;

	wire Buffer_103_clk;
	wire Buffer_103_rst;
	wire [31 : 0]Buffer_103_in1_data;
	wire Buffer_103_in1_ready;
	wire Buffer_103_in1_valid;
	wire [31 : 0]Buffer_103_out1_data;
	wire Buffer_103_out1_ready;
	wire Buffer_103_out1_valid;

	wire Buffer_104_clk;
	wire Buffer_104_rst;
	wire [31 : 0]Buffer_104_in1_data;
	wire Buffer_104_in1_ready;
	wire Buffer_104_in1_valid;
	wire [31 : 0]Buffer_104_out1_data;
	wire Buffer_104_out1_ready;
	wire Buffer_104_out1_valid;

	wire Buffer_105_clk;
	wire Buffer_105_rst;
	wire [31 : 0]Buffer_105_in1_data;
	wire Buffer_105_in1_ready;
	wire Buffer_105_in1_valid;
	wire [31 : 0]Buffer_105_out1_data;
	wire Buffer_105_out1_ready;
	wire Buffer_105_out1_valid;

	wire Buffer_106_clk;
	wire Buffer_106_rst;
	wire [31 : 0]Buffer_106_in1_data;
	wire Buffer_106_in1_ready;
	wire Buffer_106_in1_valid;
	wire [31 : 0]Buffer_106_out1_data;
	wire Buffer_106_out1_ready;
	wire Buffer_106_out1_valid;

	wire Buffer_107_clk;
	wire Buffer_107_rst;
	wire [31 : 0]Buffer_107_in1_data;
	wire Buffer_107_in1_ready;
	wire Buffer_107_in1_valid;
	wire [31 : 0]Buffer_107_out1_data;
	wire Buffer_107_out1_ready;
	wire Buffer_107_out1_valid;

	wire Buffer_108_clk;
	wire Buffer_108_rst;
	wire [31 : 0]Buffer_108_in1_data;
	wire Buffer_108_in1_ready;
	wire Buffer_108_in1_valid;
	wire [31 : 0]Buffer_108_out1_data;
	wire Buffer_108_out1_ready;
	wire Buffer_108_out1_valid;

	wire Buffer_109_clk;
	wire Buffer_109_rst;
	wire [31 : 0]Buffer_109_in1_data;
	wire Buffer_109_in1_ready;
	wire Buffer_109_in1_valid;
	wire [31 : 0]Buffer_109_out1_data;
	wire Buffer_109_out1_ready;
	wire Buffer_109_out1_valid;

	wire Buffer_110_clk;
	wire Buffer_110_rst;
	wire [31 : 0]Buffer_110_in1_data;
	wire Buffer_110_in1_ready;
	wire Buffer_110_in1_valid;
	wire [31 : 0]Buffer_110_out1_data;
	wire Buffer_110_out1_ready;
	wire Buffer_110_out1_valid;

	wire Buffer_111_clk;
	wire Buffer_111_rst;
	wire [31 : 0]Buffer_111_in1_data;
	wire Buffer_111_in1_ready;
	wire Buffer_111_in1_valid;
	wire [31 : 0]Buffer_111_out1_data;
	wire Buffer_111_out1_ready;
	wire Buffer_111_out1_valid;

	wire and_300_clk;
	wire and_300_rst;
	wire [31 : 0]and_300_in1_data;
	wire and_300_in1_ready;
	wire and_300_in1_valid;
	wire [31 : 0]and_300_in2_data;
	wire and_300_in2_ready;
	wire and_300_in2_valid;
	wire [31 : 0]and_300_out1_data;
	wire and_300_out1_ready;
	wire and_300_out1_valid;

	wire Buffer_300_clk;
	wire Buffer_300_rst;
	wire [31 : 0]Buffer_300_in1_data;
	wire Buffer_300_in1_ready;
	wire Buffer_300_in1_valid;
	wire [31 : 0]Buffer_300_out1_data;
	wire Buffer_300_out1_ready;
	wire Buffer_300_out1_valid;

	wire and_301_clk;
	wire and_301_rst;
	wire [31 : 0]and_301_in1_data;
	wire and_301_in1_ready;
	wire and_301_in1_valid;
	wire [31 : 0]and_301_in2_data;
	wire and_301_in2_ready;
	wire and_301_in2_valid;
	wire [31 : 0]and_301_out1_data;
	wire and_301_out1_ready;
	wire and_301_out1_valid;

	wire Buffer_301_clk;
	wire Buffer_301_rst;
	wire [31 : 0]Buffer_301_in1_data;
	wire Buffer_301_in1_ready;
	wire Buffer_301_in1_valid;
	wire [31 : 0]Buffer_301_out1_data;
	wire Buffer_301_out1_ready;
	wire Buffer_301_out1_valid;

	wire and_302_clk;
	wire and_302_rst;
	wire [31 : 0]and_302_in1_data;
	wire and_302_in1_ready;
	wire and_302_in1_valid;
	wire [31 : 0]and_302_in2_data;
	wire and_302_in2_ready;
	wire and_302_in2_valid;
	wire [31 : 0]and_302_out1_data;
	wire and_302_out1_ready;
	wire and_302_out1_valid;

	wire Buffer_302_clk;
	wire Buffer_302_rst;
	wire [31 : 0]Buffer_302_in1_data;
	wire Buffer_302_in1_ready;
	wire Buffer_302_in1_valid;
	wire [31 : 0]Buffer_302_out1_data;
	wire Buffer_302_out1_ready;
	wire Buffer_302_out1_valid;

	wire and_303_clk;
	wire and_303_rst;
	wire [31 : 0]and_303_in1_data;
	wire and_303_in1_ready;
	wire and_303_in1_valid;
	wire [31 : 0]and_303_in2_data;
	wire and_303_in2_ready;
	wire and_303_in2_valid;
	wire [31 : 0]and_303_out1_data;
	wire and_303_out1_ready;
	wire and_303_out1_valid;

	wire Buffer_303_clk;
	wire Buffer_303_rst;
	wire [31 : 0]Buffer_303_in1_data;
	wire Buffer_303_in1_ready;
	wire Buffer_303_in1_valid;
	wire [31 : 0]Buffer_303_out1_data;
	wire Buffer_303_out1_ready;
	wire Buffer_303_out1_valid;



	assign phi_1_clk = clk;
	assign phi_1_rst = rst;
	assign fork_0_in1_data = phi_1_out1_data;
	assign fork_0_in1_valid = phi_1_out1_valid;
	assign phi_1_out1_ready = fork_0_in1_ready;

	assign load_4_clk = clk;
	assign load_4_rst = rst;
	assign branch_1_in1_data = load_4_out1_data;
	assign branch_1_in1_valid = load_4_out1_valid;
	assign load_4_out1_ready = branch_1_in1_ready;
	assign MC_x1_in2_data = load_4_out2_data;
	assign MC_x1_in2_valid = load_4_out2_valid;
	assign load_4_out2_ready = MC_x1_in2_ready;

	assign brCst_block2_clk = clk;
	assign brCst_block2_rst = rst;
	assign fork_15_in1_data = brCst_block2_out1_data;
	assign fork_15_in1_valid = brCst_block2_out1_valid;
	assign brCst_block2_out1_ready = fork_15_in1_ready;

	assign cst_1_clk = clk;
	assign cst_1_rst = rst;
	assign branch_2_in1_data = cst_1_out1_data;
	assign branch_2_in1_valid = cst_1_out1_valid;
	assign cst_1_out1_ready = branch_2_in1_ready;

	assign fork_0_clk = clk;
	assign fork_0_rst = rst;
	assign load_4_in2_data = fork_0_out1_data;
	assign load_4_in2_valid = fork_0_out1_valid;
	assign fork_0_out1_ready = load_4_in2_ready;
	assign branch_3_in1_data = fork_0_out2_data;
	assign branch_3_in1_valid = fork_0_out2_valid;
	assign fork_0_out2_ready = branch_3_in1_ready;

	assign branch_1_clk = clk;
	assign branch_1_rst = rst;
	assign phi_6_in2_data = branch_1_out1_data;
	assign phi_6_in2_valid = branch_1_out1_valid;
	assign branch_1_out1_ready = phi_6_in2_ready;
	assign sink_1_in1_data = branch_1_out2_data;
	assign sink_1_in1_valid = branch_1_out2_valid;
	assign branch_1_out2_ready = sink_1_in1_ready;

	assign branch_2_clk = clk;
	assign branch_2_rst = rst;
	assign phi_7_in2_data = branch_2_out1_data;
	assign phi_7_in2_valid = branch_2_out1_valid;
	assign branch_2_out1_ready = phi_7_in2_ready;
	assign sink_2_in1_data = branch_2_out2_data;
	assign sink_2_in1_valid = branch_2_out2_valid;
	assign branch_2_out2_ready = sink_2_in1_ready;

	assign branch_3_clk = clk;
	assign branch_3_rst = rst;
	assign phi_n2_in1_data = branch_3_out1_data;
	assign phi_n2_in1_valid = branch_3_out1_valid;
	assign branch_3_out1_ready = phi_n2_in1_ready;
	assign sink_3_in1_data = branch_3_out2_data;
	assign sink_3_in1_valid = branch_3_out2_valid;
	assign branch_3_out2_ready = sink_3_in1_ready;

	assign fork_15_clk = clk;
	assign fork_15_rst = rst;
	assign branch_3_in2_data = fork_15_out1_data;
	assign branch_3_in2_valid = fork_15_out1_valid;
	assign fork_15_out1_ready = branch_3_in2_ready;
	assign branch_2_in2_data = fork_15_out2_data;
	assign branch_2_in2_valid = fork_15_out2_valid;
	assign fork_15_out2_ready = branch_2_in2_ready;
	assign branch_1_in2_data = fork_15_out3_data;
	assign branch_1_in2_valid = fork_15_out3_valid;
	assign fork_15_out3_ready = branch_1_in2_ready;
	assign branchC_17_in2_data = fork_15_out4_data;
	assign branchC_17_in2_valid = fork_15_out4_valid;
	assign fork_15_out4_ready = branchC_17_in2_ready;

	assign phiC_6_clk = clk;
	assign phiC_6_rst = rst;
	assign forkC_25_in1_data = phiC_6_out1_data;
	assign forkC_25_in1_valid = phiC_6_out1_valid;
	assign phiC_6_out1_ready = forkC_25_in1_ready;
	assign phi_1_in1_data = phiC_6_out2_data;
	assign phi_1_in1_valid = phiC_6_out2_valid;
	assign phiC_6_out2_ready = phi_1_in1_ready;

	assign forkC_25_clk = clk;
	assign forkC_25_rst = rst;
	assign cst_1_in1_data = forkC_25_out1_data;
	assign cst_1_in1_valid = forkC_25_out1_valid;
	assign forkC_25_out1_ready = cst_1_in1_ready;
	assign branchC_17_in1_data = forkC_25_out2_data;
	assign branchC_17_in1_valid = forkC_25_out2_valid;
	assign forkC_25_out2_ready = branchC_17_in1_ready;
	assign brCst_block2_in1_data = forkC_25_out3_data;
	assign brCst_block2_in1_valid = forkC_25_out3_valid;
	assign forkC_25_out3_ready = brCst_block2_in1_ready;

	assign branchC_17_clk = clk;
	assign branchC_17_rst = rst;
	assign phiC_7_in1_data = branchC_17_out1_data;
	assign phiC_7_in1_valid = branchC_17_out1_valid;
	assign branchC_17_out1_ready = phiC_7_in1_ready;
	assign sink_13_in1_data = branchC_17_out2_data;
	assign sink_13_in1_valid = branchC_17_out2_valid;
	assign branchC_17_out2_ready = sink_13_in1_ready;

	assign brCst_block1_clk = clk;
	assign brCst_block1_rst = rst;
	assign fork_24_in1_data = brCst_block1_out1_data;
	assign fork_24_in1_valid = brCst_block1_out1_valid;
	assign brCst_block1_out1_ready = fork_24_in1_ready;

	assign cst_0_clk = clk;
	assign cst_0_rst = rst;
	assign branch_0_in1_data = cst_0_out1_data;
	assign branch_0_in1_valid = cst_0_out1_valid;
	assign cst_0_out1_ready = branch_0_in1_ready;

	assign branch_0_clk = clk;
	assign branch_0_rst = rst;
	assign phi_1_in2_data = branch_0_out1_data;
	assign phi_1_in2_valid = branch_0_out1_valid;
	assign branch_0_out1_ready = phi_1_in2_ready;
	assign sink_0_in1_data = branch_0_out2_data;
	assign sink_0_in1_valid = branch_0_out2_valid;
	assign branch_0_out2_ready = sink_0_in1_ready;

	assign start_0_clk = clk;
	assign start_0_rst = rst;
	assign start_0_in1_data = start_in;
	assign start_0_in1_valid = start_valid;
	assign start_ready = start_0_in1_ready;
	assign forkC_23_in1_data = start_0_out1_data;
	assign forkC_23_in1_valid = start_0_out1_valid;
	assign start_0_out1_ready = forkC_23_in1_ready;

	assign forkC_23_clk = clk;
	assign forkC_23_rst = rst;
	assign cst_0_in1_data = forkC_23_out1_data;
	assign cst_0_in1_valid = forkC_23_out1_valid;
	assign forkC_23_out1_ready = cst_0_in1_ready;
	assign branchC_16_in1_data = forkC_23_out2_data;
	assign branchC_16_in1_valid = forkC_23_out2_valid;
	assign forkC_23_out2_ready = branchC_16_in1_ready;
	assign brCst_block1_in1_data = forkC_23_out3_data;
	assign brCst_block1_in1_valid = forkC_23_out3_valid;
	assign forkC_23_out3_ready = brCst_block1_in1_ready;

	assign branchC_16_clk = clk;
	assign branchC_16_rst = rst;
	assign phiC_6_in1_data = branchC_16_out1_data;
	assign phiC_6_in1_valid = branchC_16_out1_valid;
	assign branchC_16_out1_ready = phiC_6_in1_ready;
	assign sink_12_in1_data = branchC_16_out2_data;
	assign sink_12_in1_valid = branchC_16_out2_valid;
	assign branchC_16_out2_ready = sink_12_in1_ready;

	assign fork_24_clk = clk;
	assign fork_24_rst = rst;
	assign branch_0_in2_data = fork_24_out1_data;
	assign branch_0_in2_valid = fork_24_out1_valid;
	assign fork_24_out1_ready = branch_0_in2_ready;
	assign branchC_16_in2_data = fork_24_out2_data;
	assign branchC_16_in2_valid = fork_24_out2_valid;
	assign fork_24_out2_ready = branchC_16_in2_ready;

	assign phi_27_clk = clk;
	assign phi_27_rst = rst;
	assign fork_5_in1_data = phi_27_out1_data;
	assign fork_5_in1_valid = phi_27_out1_valid;
	assign phi_27_out1_ready = fork_5_in1_ready;

	assign load_30_clk = clk;
	assign load_30_rst = rst;
	assign branch_9_in1_data = load_30_out1_data;
	assign branch_9_in1_valid = load_30_out1_valid;
	assign load_30_out1_ready = branch_9_in1_ready;
	assign MC_x2_in2_data = load_30_out2_data;
	assign MC_x2_in2_valid = load_30_out2_valid;
	assign load_30_out2_ready = MC_x2_in2_ready;

	assign brCst_block6_clk = clk;
	assign brCst_block6_rst = rst;
	assign fork_19_in1_data = brCst_block6_out1_data;
	assign fork_19_in1_valid = brCst_block6_out1_valid;
	assign brCst_block6_out1_ready = fork_19_in1_ready;

	assign cst_8_clk = clk;
	assign cst_8_rst = rst;
	assign branch_10_in1_data = cst_8_out1_data;
	assign branch_10_in1_valid = cst_8_out1_valid;
	assign cst_8_out1_ready = branch_10_in1_ready;

	assign fork_5_clk = clk;
	assign fork_5_rst = rst;
	assign load_30_in2_data = fork_5_out1_data;
	assign load_30_in2_valid = fork_5_out1_valid;
	assign fork_5_out1_ready = load_30_in2_ready;
	assign branch_11_in1_data = fork_5_out2_data;
	assign branch_11_in1_valid = fork_5_out2_valid;
	assign fork_5_out2_ready = branch_11_in1_ready;

	assign branch_9_clk = clk;
	assign branch_9_rst = rst;
	assign phi_32_in2_data = branch_9_out1_data;
	assign phi_32_in2_valid = branch_9_out1_valid;
	assign branch_9_out1_ready = phi_32_in2_ready;
	assign sink_7_in1_data = branch_9_out2_data;
	assign sink_7_in1_valid = branch_9_out2_valid;
	assign branch_9_out2_ready = sink_7_in1_ready;

	assign branch_10_clk = clk;
	assign branch_10_rst = rst;
	assign phi_33_in2_data = branch_10_out1_data;
	assign phi_33_in2_valid = branch_10_out1_valid;
	assign branch_10_out1_ready = phi_33_in2_ready;
	assign sink_8_in1_data = branch_10_out2_data;
	assign sink_8_in1_valid = branch_10_out2_valid;
	assign branch_10_out2_ready = sink_8_in1_ready;

	assign branch_11_clk = clk;
	assign branch_11_rst = rst;
	assign phi_n5_in1_data = branch_11_out1_data;
	assign phi_n5_in1_valid = branch_11_out1_valid;
	assign branch_11_out1_ready = phi_n5_in1_ready;
	assign sink_9_in1_data = branch_11_out2_data;
	assign sink_9_in1_valid = branch_11_out2_valid;
	assign branch_11_out2_ready = sink_9_in1_ready;

	assign fork_19_clk = clk;
	assign fork_19_rst = rst;
	assign branch_11_in2_data = fork_19_out1_data;
	assign branch_11_in2_valid = fork_19_out1_valid;
	assign fork_19_out1_ready = branch_11_in2_ready;
	assign branch_10_in2_data = fork_19_out2_data;
	assign branch_10_in2_valid = fork_19_out2_valid;
	assign fork_19_out2_ready = branch_10_in2_ready;
	assign branch_9_in2_data = fork_19_out3_data;
	assign branch_9_in2_valid = fork_19_out3_valid;
	assign fork_19_out3_ready = branch_9_in2_ready;
	assign branchC_21_in2_data = fork_19_out4_data;
	assign branchC_21_in2_valid = fork_19_out4_valid;
	assign fork_19_out4_ready = branchC_21_in2_ready;

	assign phiC_10_clk = clk;
	assign phiC_10_rst = rst;
	assign forkC_31_in1_data = phiC_10_out1_data;
	assign forkC_31_in1_valid = phiC_10_out1_valid;
	assign phiC_10_out1_ready = forkC_31_in1_ready;
	assign phi_27_in1_data = phiC_10_out2_data;
	assign phi_27_in1_valid = phiC_10_out2_valid;
	assign phiC_10_out2_ready = phi_27_in1_ready;

	assign forkC_31_clk = clk;
	assign forkC_31_rst = rst;
	assign cst_8_in1_data = forkC_31_out1_data;
	assign cst_8_in1_valid = forkC_31_out1_valid;
	assign forkC_31_out1_ready = cst_8_in1_ready;
	assign branchC_21_in1_data = forkC_31_out2_data;
	assign branchC_21_in1_valid = forkC_31_out2_valid;
	assign forkC_31_out2_ready = branchC_21_in1_ready;
	assign brCst_block6_in1_data = forkC_31_out3_data;
	assign brCst_block6_in1_valid = forkC_31_out3_valid;
	assign forkC_31_out3_ready = brCst_block6_in1_ready;

	assign branchC_21_clk = clk;
	assign branchC_21_rst = rst;
	assign phiC_11_in1_data = branchC_21_out1_data;
	assign phiC_11_in1_valid = branchC_21_out1_valid;
	assign branchC_21_out1_ready = phiC_11_in1_ready;
	assign sink_15_in1_data = branchC_21_out2_data;
	assign sink_15_in1_valid = branchC_21_out2_valid;
	assign branchC_21_out2_ready = sink_15_in1_ready;

	assign phi_32_clk = clk;
	assign phi_32_rst = rst;
	assign and_303_in1_data = phi_32_out1_data;
	assign and_303_in1_valid = phi_32_out1_valid;
	assign phi_32_out1_ready = and_303_in1_ready;

	assign phi_33_clk = clk;
	assign phi_33_rst = rst;
	assign fork_6_in1_data = phi_33_out1_data;
	assign fork_6_in1_valid = phi_33_out1_valid;
	assign phi_33_out1_ready = fork_6_in1_ready;

	assign cst_9_clk = clk;
	assign cst_9_rst = rst;
	assign shl_34_in2_data = cst_9_out1_data;
	assign shl_34_in2_valid = cst_9_out1_valid;
	assign cst_9_out1_ready = shl_34_in2_ready;

	assign shl_34_clk = clk;
	assign shl_34_rst = rst;
	assign add_35_in1_data = shl_34_out1_data;
	assign add_35_in1_valid = shl_34_out1_valid;
	assign shl_34_out1_ready = add_35_in1_ready;

	assign add_35_clk = clk;
	assign add_35_rst = rst;
	assign load_38_in2_data = add_35_out1_data;
	assign load_38_in2_valid = add_35_out1_valid;
	assign add_35_out1_ready = load_38_in2_ready;

	assign load_38_clk = clk;
	assign load_38_rst = rst;
	assign and_302_in1_data = load_38_out1_data;
	assign and_302_in1_valid = load_38_out1_valid;
	assign load_38_out1_ready = and_302_in1_ready;
	assign MC_A_in2_data = load_38_out2_data;
	assign MC_A_in2_valid = load_38_out2_valid;
	assign load_38_out2_ready = MC_A_in2_ready;

	assign load_41_clk = clk;
	assign load_41_rst = rst;
	assign and_302_in2_data = load_41_out1_data;
	assign and_302_in2_valid = load_41_out1_valid;
	assign load_41_out1_ready = and_302_in2_ready;
	assign MC_y2_in1_data = load_41_out2_data;
	assign MC_y2_in1_valid = load_41_out2_valid;
	assign load_41_out2_ready = MC_y2_in1_ready;

	assign cst_10_clk = clk;
	assign cst_10_rst = rst;
	assign add_44_in2_data = cst_10_out1_data;
	assign add_44_in2_valid = cst_10_out1_valid;
	assign cst_10_out1_ready = add_44_in2_ready;

	assign add_44_clk = clk;
	assign add_44_rst = rst;
	assign fork_8_in1_data = add_44_out1_data;
	assign fork_8_in1_valid = add_44_out1_valid;
	assign add_44_out1_ready = fork_8_in1_ready;

	assign cst_11_clk = clk;
	assign cst_11_rst = rst;
	assign icmp_45_in2_data = cst_11_out1_data;
	assign icmp_45_in2_valid = cst_11_out1_valid;
	assign cst_11_out1_ready = icmp_45_in2_ready;

	assign icmp_45_clk = clk;
	assign icmp_45_rst = rst;
	assign fork_20_in1_data = icmp_45_out1_data;
	assign fork_20_in1_valid = icmp_45_out1_valid;
	assign icmp_45_out1_ready = fork_20_in1_ready;

	assign phi_n5_clk = clk;
	assign phi_n5_rst = rst;
	assign fork_13_in1_data = phi_n5_out1_data;
	assign fork_13_in1_valid = phi_n5_out1_valid;
	assign phi_n5_out1_ready = fork_13_in1_ready;

	assign fork_6_clk = clk;
	assign fork_6_rst = rst;
	assign shl_34_in1_data = fork_6_out1_data;
	assign shl_34_in1_valid = fork_6_out1_valid;
	assign fork_6_out1_ready = shl_34_in1_ready;
	assign add_44_in1_data = fork_6_out2_data;
	assign add_44_in1_valid = fork_6_out2_valid;
	assign fork_6_out2_ready = add_44_in1_ready;
	assign load_41_in2_data = fork_6_out3_data;
	assign load_41_in2_valid = fork_6_out3_valid;
	assign fork_6_out3_ready = load_41_in2_ready;

	assign fork_8_clk = clk;
	assign fork_8_rst = rst;
	assign icmp_45_in1_data = fork_8_out1_data;
	assign icmp_45_in1_valid = fork_8_out1_valid;
	assign fork_8_out1_ready = icmp_45_in1_ready;
	assign branch_13_in1_data = fork_8_out2_data;
	assign branch_13_in1_valid = fork_8_out2_valid;
	assign fork_8_out2_ready = branch_13_in1_ready;

	assign fork_13_clk = clk;
	assign fork_13_rst = rst;
	assign add_35_in2_data = fork_13_out1_data;
	assign add_35_in2_valid = fork_13_out1_valid;
	assign fork_13_out1_ready = add_35_in2_ready;
	assign branch_14_in1_data = fork_13_out2_data;
	assign branch_14_in1_valid = fork_13_out2_valid;
	assign fork_13_out2_ready = branch_14_in1_ready;

	assign branch_12_clk = clk;
	assign branch_12_rst = rst;
	assign Buffer_106_in1_data = branch_12_out1_data;
	assign Buffer_106_in1_valid = branch_12_out1_valid;
	assign branch_12_out1_ready = Buffer_106_in1_ready;
	assign phi_n3_in1_data = branch_12_out2_data;
	assign phi_n3_in1_valid = branch_12_out2_valid;
	assign branch_12_out2_ready = phi_n3_in1_ready;

	assign branch_13_clk = clk;
	assign branch_13_rst = rst;
	assign Buffer_107_in1_data = branch_13_out1_data;
	assign Buffer_107_in1_valid = branch_13_out1_valid;
	assign branch_13_out1_ready = Buffer_107_in1_ready;
	assign sink_10_in1_data = branch_13_out2_data;
	assign sink_10_in1_valid = branch_13_out2_valid;
	assign branch_13_out2_ready = sink_10_in1_ready;

	assign branch_14_clk = clk;
	assign branch_14_rst = rst;
	assign Buffer_108_in1_data = branch_14_out1_data;
	assign Buffer_108_in1_valid = branch_14_out1_valid;
	assign branch_14_out1_ready = Buffer_108_in1_ready;
	assign phi_n4_in1_data = branch_14_out2_data;
	assign phi_n4_in1_valid = branch_14_out2_valid;
	assign branch_14_out2_ready = phi_n4_in1_ready;

	assign fork_20_clk = clk;
	assign fork_20_rst = rst;
	assign branch_14_in2_data = fork_20_out1_data;
	assign branch_14_in2_valid = fork_20_out1_valid;
	assign fork_20_out1_ready = branch_14_in2_ready;
	assign branch_13_in2_data = fork_20_out2_data;
	assign branch_13_in2_valid = fork_20_out2_valid;
	assign fork_20_out2_ready = branch_13_in2_ready;
	assign branch_12_in2_data = fork_20_out3_data;
	assign branch_12_in2_valid = fork_20_out3_valid;
	assign fork_20_out3_ready = branch_12_in2_ready;
	assign branchC_22_in2_data = fork_20_out4_data;
	assign branchC_22_in2_valid = fork_20_out4_valid;
	assign fork_20_out4_ready = branchC_22_in2_ready;

	assign phiC_11_clk = clk;
	assign phiC_11_rst = rst;
	assign branchC_22_in1_data = phiC_11_out1_data;
	assign branchC_22_in1_valid = phiC_11_out1_valid;
	assign phiC_11_out1_ready = branchC_22_in1_ready;
	assign fork_39_in1_data = phiC_11_out2_data;
	assign fork_39_in1_valid = phiC_11_out2_valid;
	assign phiC_11_out2_ready = fork_39_in1_ready;

	assign branchC_22_clk = clk;
	assign branchC_22_rst = rst;
	assign Buffer_109_in1_data = branchC_22_out1_data;
	assign Buffer_109_in1_valid = branchC_22_out1_valid;
	assign branchC_22_out1_ready = Buffer_109_in1_ready;
	assign phiC_12_in1_data = branchC_22_out2_data;
	assign phiC_12_in1_valid = branchC_22_out2_valid;
	assign branchC_22_out2_ready = phiC_12_in1_ready;

	assign source_5_clk = clk;
	assign source_5_rst = rst;
	assign cst_9_in1_data = source_5_out1_data;
	assign cst_9_in1_valid = source_5_out1_valid;
	assign source_5_out1_ready = cst_9_in1_ready;

	assign source_6_clk = clk;
	assign source_6_rst = rst;
	assign cst_10_in1_data = source_6_out1_data;
	assign cst_10_in1_valid = source_6_out1_valid;
	assign source_6_out1_ready = cst_10_in1_ready;

	assign source_7_clk = clk;
	assign source_7_rst = rst;
	assign cst_11_in1_data = source_7_out1_data;
	assign cst_11_in1_valid = source_7_out1_valid;
	assign source_7_out1_ready = cst_11_in1_ready;

	assign fork_39_clk = clk;
	assign fork_39_rst = rst;
	assign phi_32_in1_data = fork_39_out1_data;
	assign phi_32_in1_valid = fork_39_out1_valid;
	assign fork_39_out1_ready = phi_32_in1_ready;
	assign phi_33_in1_data = fork_39_out2_data;
	assign phi_33_in1_valid = fork_39_out2_valid;
	assign fork_39_out2_ready = phi_33_in1_ready;

	assign store_1_clk = clk;
	assign store_1_rst = rst;
	assign MC_x2_in4_data = store_1_out1_data;
	assign MC_x2_in4_valid = store_1_out1_valid;
	assign store_1_out1_ready = MC_x2_in4_ready;
	assign MC_x2_in3_data = store_1_out2_data;
	assign MC_x2_in3_valid = store_1_out2_valid;
	assign store_1_out2_ready = MC_x2_in3_ready;

	assign cst_12_clk = clk;
	assign cst_12_rst = rst;
	assign add_49_in2_data = cst_12_out1_data;
	assign add_49_in2_valid = cst_12_out1_valid;
	assign cst_12_out1_ready = add_49_in2_ready;

	assign add_49_clk = clk;
	assign add_49_rst = rst;
	assign fork_9_in1_data = add_49_out1_data;
	assign fork_9_in1_valid = add_49_out1_valid;
	assign add_49_out1_ready = fork_9_in1_ready;

	assign cst_13_clk = clk;
	assign cst_13_rst = rst;
	assign icmp_50_in2_data = cst_13_out1_data;
	assign icmp_50_in2_valid = cst_13_out1_valid;
	assign cst_13_out1_ready = icmp_50_in2_ready;

	assign icmp_50_clk = clk;
	assign icmp_50_rst = rst;
	assign fork_34_in1_data = icmp_50_out1_data;
	assign fork_34_in1_valid = icmp_50_out1_valid;
	assign icmp_50_out1_ready = fork_34_in1_ready;

	assign phi_n3_clk = clk;
	assign phi_n3_rst = rst;
	assign store_1_in1_data = phi_n3_out1_data;
	assign store_1_in1_valid = phi_n3_out1_valid;
	assign phi_n3_out1_ready = store_1_in1_ready;

	assign phi_n4_clk = clk;
	assign phi_n4_rst = rst;
	assign fork_12_in1_data = phi_n4_out1_data;
	assign fork_12_in1_valid = phi_n4_out1_valid;
	assign phi_n4_out1_ready = fork_12_in1_ready;

	assign fork_9_clk = clk;
	assign fork_9_rst = rst;
	assign icmp_50_in1_data = fork_9_out1_data;
	assign icmp_50_in1_valid = fork_9_out1_valid;
	assign fork_9_out1_ready = icmp_50_in1_ready;
	assign branch_15_in1_data = fork_9_out2_data;
	assign branch_15_in1_valid = fork_9_out2_valid;
	assign fork_9_out2_ready = branch_15_in1_ready;

	assign fork_12_clk = clk;
	assign fork_12_rst = rst;
	assign store_1_in2_data = fork_12_out1_data;
	assign store_1_in2_valid = fork_12_out1_valid;
	assign fork_12_out1_ready = store_1_in2_ready;
	assign add_49_in1_data = fork_12_out2_data;
	assign add_49_in1_valid = fork_12_out2_valid;
	assign fork_12_out2_ready = add_49_in1_ready;

	assign branch_15_clk = clk;
	assign branch_15_rst = rst;
	assign Buffer_110_in1_data = branch_15_out1_data;
	assign Buffer_110_in1_valid = branch_15_out1_valid;
	assign branch_15_out1_ready = Buffer_110_in1_ready;
	assign sink_11_in1_data = branch_15_out2_data;
	assign sink_11_in1_valid = branch_15_out2_valid;
	assign branch_15_out2_ready = sink_11_in1_ready;

	assign cst_15_clk = clk;
	assign cst_15_rst = rst;
	assign MC_x2_in1_data = cst_15_out1_data;
	assign MC_x2_in1_valid = cst_15_out1_valid;
	assign cst_15_out1_ready = MC_x2_in1_ready;

	assign phiC_12_clk = clk;
	assign phiC_12_rst = rst;
	assign forkC_33_in1_data = phiC_12_out1_data;
	assign forkC_33_in1_valid = phiC_12_out1_valid;
	assign phiC_12_out1_ready = forkC_33_in1_ready;

	assign forkC_33_clk = clk;
	assign forkC_33_rst = rst;
	assign cst_15_in1_data = forkC_33_out1_data;
	assign cst_15_in1_valid = forkC_33_out1_valid;
	assign forkC_33_out1_ready = cst_15_in1_ready;
	assign branchC_23_in1_data = forkC_33_out2_data;
	assign branchC_23_in1_valid = forkC_33_out2_valid;
	assign forkC_33_out2_ready = branchC_23_in1_ready;

	assign branchC_23_clk = clk;
	assign branchC_23_rst = rst;
	assign Buffer_111_in1_data = branchC_23_out1_data;
	assign Buffer_111_in1_valid = branchC_23_out1_valid;
	assign branchC_23_out1_ready = Buffer_111_in1_ready;
	assign phiC_13_in1_data = branchC_23_out2_data;
	assign phiC_13_in1_valid = branchC_23_out2_valid;
	assign branchC_23_out2_ready = phiC_13_in1_ready;

	assign fork_34_clk = clk;
	assign fork_34_rst = rst;
	assign branch_15_in2_data = fork_34_out1_data;
	assign branch_15_in2_valid = fork_34_out1_valid;
	assign fork_34_out1_ready = branch_15_in2_ready;
	assign branchC_23_in2_data = fork_34_out2_data;
	assign branchC_23_in2_valid = fork_34_out2_valid;
	assign fork_34_out2_ready = branchC_23_in2_ready;

	assign source_8_clk = clk;
	assign source_8_rst = rst;
	assign cst_12_in1_data = source_8_out1_data;
	assign cst_12_in1_valid = source_8_out1_valid;
	assign source_8_out1_ready = cst_12_in1_ready;

	assign source_9_clk = clk;
	assign source_9_rst = rst;
	assign cst_13_in1_data = source_9_out1_data;
	assign cst_13_in1_valid = source_9_out1_valid;
	assign source_9_out1_ready = cst_13_in1_ready;

	assign brCst_block5_clk = clk;
	assign brCst_block5_rst = rst;
	assign fork_30_in1_data = brCst_block5_out1_data;
	assign fork_30_in1_valid = brCst_block5_out1_valid;
	assign brCst_block5_out1_ready = fork_30_in1_ready;

	assign cst_7_clk = clk;
	assign cst_7_rst = rst;
	assign branch_8_in1_data = cst_7_out1_data;
	assign branch_8_in1_valid = cst_7_out1_valid;
	assign cst_7_out1_ready = branch_8_in1_ready;

	assign branch_8_clk = clk;
	assign branch_8_rst = rst;
	assign phi_27_in2_data = branch_8_out1_data;
	assign phi_27_in2_valid = branch_8_out1_valid;
	assign branch_8_out1_ready = phi_27_in2_ready;
	assign sink_6_in1_data = branch_8_out2_data;
	assign sink_6_in1_valid = branch_8_out2_valid;
	assign branch_8_out2_ready = sink_6_in1_ready;

	assign phiC_9_clk = clk;
	assign phiC_9_rst = rst;
	assign forkC_29_in1_data = phiC_9_out1_data;
	assign forkC_29_in1_valid = phiC_9_out1_valid;
	assign phiC_9_out1_ready = forkC_29_in1_ready;

	assign forkC_29_clk = clk;
	assign forkC_29_rst = rst;
	assign cst_7_in1_data = forkC_29_out1_data;
	assign cst_7_in1_valid = forkC_29_out1_valid;
	assign forkC_29_out1_ready = cst_7_in1_ready;
	assign branchC_20_in1_data = forkC_29_out2_data;
	assign branchC_20_in1_valid = forkC_29_out2_valid;
	assign forkC_29_out2_ready = branchC_20_in1_ready;
	assign brCst_block5_in1_data = forkC_29_out3_data;
	assign brCst_block5_in1_valid = forkC_29_out3_valid;
	assign forkC_29_out3_ready = brCst_block5_in1_ready;

	assign branchC_20_clk = clk;
	assign branchC_20_rst = rst;
	assign phiC_10_in1_data = branchC_20_out1_data;
	assign phiC_10_in1_valid = branchC_20_out1_valid;
	assign branchC_20_out1_ready = phiC_10_in1_ready;
	assign sink_14_in1_data = branchC_20_out2_data;
	assign sink_14_in1_valid = branchC_20_out2_valid;
	assign branchC_20_out2_ready = sink_14_in1_ready;

	assign fork_30_clk = clk;
	assign fork_30_rst = rst;
	assign branch_8_in2_data = fork_30_out1_data;
	assign branch_8_in2_valid = fork_30_out1_valid;
	assign fork_30_out1_ready = branch_8_in2_ready;
	assign branchC_20_in2_data = fork_30_out2_data;
	assign branchC_20_in2_valid = fork_30_out2_valid;
	assign fork_30_out2_ready = branchC_20_in2_ready;

	assign phi_6_clk = clk;
	assign phi_6_rst = rst;
	assign and_301_in1_data = phi_6_out1_data;
	assign and_301_in1_valid = phi_6_out1_valid;
	assign phi_6_out1_ready = and_301_in1_ready;

	assign phi_7_clk = clk;
	assign phi_7_rst = rst;
	assign fork_1_in1_data = phi_7_out1_data;
	assign fork_1_in1_valid = phi_7_out1_valid;
	assign phi_7_out1_ready = fork_1_in1_ready;

	assign cst_2_clk = clk;
	assign cst_2_rst = rst;
	assign shl_8_in2_data = cst_2_out1_data;
	assign shl_8_in2_valid = cst_2_out1_valid;
	assign cst_2_out1_ready = shl_8_in2_ready;

	assign shl_8_clk = clk;
	assign shl_8_rst = rst;
	assign add_9_in1_data = shl_8_out1_data;
	assign add_9_in1_valid = shl_8_out1_valid;
	assign shl_8_out1_ready = add_9_in1_ready;

	assign add_9_clk = clk;
	assign add_9_rst = rst;
	assign load_12_in2_data = add_9_out1_data;
	assign load_12_in2_valid = add_9_out1_valid;
	assign add_9_out1_ready = load_12_in2_ready;

	assign load_12_clk = clk;
	assign load_12_rst = rst;
	assign and_300_in1_data = load_12_out1_data;
	assign and_300_in1_valid = load_12_out1_valid;
	assign load_12_out1_ready = and_300_in1_ready;
	assign MC_A_in1_data = load_12_out2_data;
	assign MC_A_in1_valid = load_12_out2_valid;
	assign load_12_out2_ready = MC_A_in1_ready;

	assign load_15_clk = clk;
	assign load_15_rst = rst;
	assign and_300_in2_data = load_15_out1_data;
	assign and_300_in2_valid = load_15_out1_valid;
	assign load_15_out1_ready = and_300_in2_ready;
	assign MC_y1_in1_data = load_15_out2_data;
	assign MC_y1_in1_valid = load_15_out2_valid;
	assign load_15_out2_ready = MC_y1_in1_ready;

	assign cst_3_clk = clk;
	assign cst_3_rst = rst;
	assign add_18_in2_data = cst_3_out1_data;
	assign add_18_in2_valid = cst_3_out1_valid;
	assign cst_3_out1_ready = add_18_in2_ready;

	assign add_18_clk = clk;
	assign add_18_rst = rst;
	assign fork_3_in1_data = add_18_out1_data;
	assign fork_3_in1_valid = add_18_out1_valid;
	assign add_18_out1_ready = fork_3_in1_ready;

	assign cst_4_clk = clk;
	assign cst_4_rst = rst;
	assign icmp_19_in2_data = cst_4_out1_data;
	assign icmp_19_in2_valid = cst_4_out1_valid;
	assign cst_4_out1_ready = icmp_19_in2_ready;

	assign icmp_19_clk = clk;
	assign icmp_19_rst = rst;
	assign fork_16_in1_data = icmp_19_out1_data;
	assign fork_16_in1_valid = icmp_19_out1_valid;
	assign icmp_19_out1_ready = fork_16_in1_ready;

	assign phi_n2_clk = clk;
	assign phi_n2_rst = rst;
	assign fork_11_in1_data = phi_n2_out1_data;
	assign fork_11_in1_valid = phi_n2_out1_valid;
	assign phi_n2_out1_ready = fork_11_in1_ready;

	assign fork_1_clk = clk;
	assign fork_1_rst = rst;
	assign add_9_in2_data = fork_1_out1_data;
	assign add_9_in2_valid = fork_1_out1_valid;
	assign fork_1_out1_ready = add_9_in2_ready;
	assign add_18_in1_data = fork_1_out2_data;
	assign add_18_in1_valid = fork_1_out2_valid;
	assign fork_1_out2_ready = add_18_in1_ready;
	assign load_15_in2_data = fork_1_out3_data;
	assign load_15_in2_valid = fork_1_out3_valid;
	assign fork_1_out3_ready = load_15_in2_ready;

	assign fork_3_clk = clk;
	assign fork_3_rst = rst;
	assign icmp_19_in1_data = fork_3_out1_data;
	assign icmp_19_in1_valid = fork_3_out1_valid;
	assign fork_3_out1_ready = icmp_19_in1_ready;
	assign branch_5_in1_data = fork_3_out2_data;
	assign branch_5_in1_valid = fork_3_out2_valid;
	assign fork_3_out2_ready = branch_5_in1_ready;

	assign fork_11_clk = clk;
	assign fork_11_rst = rst;
	assign shl_8_in1_data = fork_11_out1_data;
	assign shl_8_in1_valid = fork_11_out1_valid;
	assign fork_11_out1_ready = shl_8_in1_ready;
	assign branch_6_in1_data = fork_11_out2_data;
	assign branch_6_in1_valid = fork_11_out2_valid;
	assign fork_11_out2_ready = branch_6_in1_ready;

	assign branch_4_clk = clk;
	assign branch_4_rst = rst;
	assign Buffer_100_in1_data = branch_4_out1_data;
	assign Buffer_100_in1_valid = branch_4_out1_valid;
	assign branch_4_out1_ready = Buffer_100_in1_ready;
	assign phi_n0_in1_data = branch_4_out2_data;
	assign phi_n0_in1_valid = branch_4_out2_valid;
	assign branch_4_out2_ready = phi_n0_in1_ready;

	assign branch_5_clk = clk;
	assign branch_5_rst = rst;
	assign Buffer_101_in1_data = branch_5_out1_data;
	assign Buffer_101_in1_valid = branch_5_out1_valid;
	assign branch_5_out1_ready = Buffer_101_in1_ready;
	assign sink_4_in1_data = branch_5_out2_data;
	assign sink_4_in1_valid = branch_5_out2_valid;
	assign branch_5_out2_ready = sink_4_in1_ready;

	assign branch_6_clk = clk;
	assign branch_6_rst = rst;
	assign Buffer_102_in1_data = branch_6_out1_data;
	assign Buffer_102_in1_valid = branch_6_out1_valid;
	assign branch_6_out1_ready = Buffer_102_in1_ready;
	assign phi_n1_in1_data = branch_6_out2_data;
	assign phi_n1_in1_valid = branch_6_out2_valid;
	assign branch_6_out2_ready = phi_n1_in1_ready;

	assign fork_16_clk = clk;
	assign fork_16_rst = rst;
	assign branch_6_in2_data = fork_16_out1_data;
	assign branch_6_in2_valid = fork_16_out1_valid;
	assign fork_16_out1_ready = branch_6_in2_ready;
	assign branch_5_in2_data = fork_16_out2_data;
	assign branch_5_in2_valid = fork_16_out2_valid;
	assign fork_16_out2_ready = branch_5_in2_ready;
	assign branch_4_in2_data = fork_16_out3_data;
	assign branch_4_in2_valid = fork_16_out3_valid;
	assign fork_16_out3_ready = branch_4_in2_ready;
	assign branchC_18_in2_data = fork_16_out4_data;
	assign branchC_18_in2_valid = fork_16_out4_valid;
	assign fork_16_out4_ready = branchC_18_in2_ready;

	assign phiC_7_clk = clk;
	assign phiC_7_rst = rst;
	assign branchC_18_in1_data = phiC_7_out1_data;
	assign branchC_18_in1_valid = phiC_7_out1_valid;
	assign phiC_7_out1_ready = branchC_18_in1_ready;
	assign fork_37_in1_data = phiC_7_out2_data;
	assign fork_37_in1_valid = phiC_7_out2_valid;
	assign phiC_7_out2_ready = fork_37_in1_ready;

	assign branchC_18_clk = clk;
	assign branchC_18_rst = rst;
	assign Buffer_103_in1_data = branchC_18_out1_data;
	assign Buffer_103_in1_valid = branchC_18_out1_valid;
	assign branchC_18_out1_ready = Buffer_103_in1_ready;
	assign phiC_8_in1_data = branchC_18_out2_data;
	assign phiC_8_in1_valid = branchC_18_out2_valid;
	assign branchC_18_out2_ready = phiC_8_in1_ready;

	assign source_0_clk = clk;
	assign source_0_rst = rst;
	assign cst_2_in1_data = source_0_out1_data;
	assign cst_2_in1_valid = source_0_out1_valid;
	assign source_0_out1_ready = cst_2_in1_ready;

	assign source_1_clk = clk;
	assign source_1_rst = rst;
	assign cst_3_in1_data = source_1_out1_data;
	assign cst_3_in1_valid = source_1_out1_valid;
	assign source_1_out1_ready = cst_3_in1_ready;

	assign source_2_clk = clk;
	assign source_2_rst = rst;
	assign cst_4_in1_data = source_2_out1_data;
	assign cst_4_in1_valid = source_2_out1_valid;
	assign source_2_out1_ready = cst_4_in1_ready;

	assign fork_37_clk = clk;
	assign fork_37_rst = rst;
	assign phi_6_in1_data = fork_37_out1_data;
	assign phi_6_in1_valid = fork_37_out1_valid;
	assign fork_37_out1_ready = phi_6_in1_ready;
	assign phi_7_in1_data = fork_37_out2_data;
	assign phi_7_in1_valid = fork_37_out2_valid;
	assign fork_37_out2_ready = phi_7_in1_ready;

	assign store_0_clk = clk;
	assign store_0_rst = rst;
	assign MC_x1_in4_data = store_0_out1_data;
	assign MC_x1_in4_valid = store_0_out1_valid;
	assign store_0_out1_ready = MC_x1_in4_ready;
	assign MC_x1_in3_data = store_0_out2_data;
	assign MC_x1_in3_valid = store_0_out2_valid;
	assign store_0_out2_ready = MC_x1_in3_ready;

	assign cst_5_clk = clk;
	assign cst_5_rst = rst;
	assign add_23_in2_data = cst_5_out1_data;
	assign add_23_in2_valid = cst_5_out1_valid;
	assign cst_5_out1_ready = add_23_in2_ready;

	assign add_23_clk = clk;
	assign add_23_rst = rst;
	assign fork_4_in1_data = add_23_out1_data;
	assign fork_4_in1_valid = add_23_out1_valid;
	assign add_23_out1_ready = fork_4_in1_ready;

	assign cst_6_clk = clk;
	assign cst_6_rst = rst;
	assign icmp_24_in2_data = cst_6_out1_data;
	assign icmp_24_in2_valid = cst_6_out1_valid;
	assign cst_6_out1_ready = icmp_24_in2_ready;

	assign icmp_24_clk = clk;
	assign icmp_24_rst = rst;
	assign fork_28_in1_data = icmp_24_out1_data;
	assign fork_28_in1_valid = icmp_24_out1_valid;
	assign icmp_24_out1_ready = fork_28_in1_ready;

	assign phi_n0_clk = clk;
	assign phi_n0_rst = rst;
	assign store_0_in1_data = phi_n0_out1_data;
	assign store_0_in1_valid = phi_n0_out1_valid;
	assign phi_n0_out1_ready = store_0_in1_ready;

	assign phi_n1_clk = clk;
	assign phi_n1_rst = rst;
	assign fork_10_in1_data = phi_n1_out1_data;
	assign fork_10_in1_valid = phi_n1_out1_valid;
	assign phi_n1_out1_ready = fork_10_in1_ready;

	assign fork_4_clk = clk;
	assign fork_4_rst = rst;
	assign icmp_24_in1_data = fork_4_out1_data;
	assign icmp_24_in1_valid = fork_4_out1_valid;
	assign fork_4_out1_ready = icmp_24_in1_ready;
	assign branch_7_in1_data = fork_4_out2_data;
	assign branch_7_in1_valid = fork_4_out2_valid;
	assign fork_4_out2_ready = branch_7_in1_ready;

	assign fork_10_clk = clk;
	assign fork_10_rst = rst;
	assign store_0_in2_data = fork_10_out1_data;
	assign store_0_in2_valid = fork_10_out1_valid;
	assign fork_10_out1_ready = store_0_in2_ready;
	assign add_23_in1_data = fork_10_out2_data;
	assign add_23_in1_valid = fork_10_out2_valid;
	assign fork_10_out2_ready = add_23_in1_ready;

	assign branch_7_clk = clk;
	assign branch_7_rst = rst;
	assign Buffer_104_in1_data = branch_7_out1_data;
	assign Buffer_104_in1_valid = branch_7_out1_valid;
	assign branch_7_out1_ready = Buffer_104_in1_ready;
	assign sink_5_in1_data = branch_7_out2_data;
	assign sink_5_in1_valid = branch_7_out2_valid;
	assign branch_7_out2_ready = sink_5_in1_ready;

	assign cst_14_clk = clk;
	assign cst_14_rst = rst;
	assign MC_x1_in1_data = cst_14_out1_data;
	assign MC_x1_in1_valid = cst_14_out1_valid;
	assign cst_14_out1_ready = MC_x1_in1_ready;

	assign phiC_8_clk = clk;
	assign phiC_8_rst = rst;
	assign forkC_27_in1_data = phiC_8_out1_data;
	assign forkC_27_in1_valid = phiC_8_out1_valid;
	assign phiC_8_out1_ready = forkC_27_in1_ready;

	assign forkC_27_clk = clk;
	assign forkC_27_rst = rst;
	assign cst_14_in1_data = forkC_27_out1_data;
	assign cst_14_in1_valid = forkC_27_out1_valid;
	assign forkC_27_out1_ready = cst_14_in1_ready;
	assign branchC_19_in1_data = forkC_27_out2_data;
	assign branchC_19_in1_valid = forkC_27_out2_valid;
	assign forkC_27_out2_ready = branchC_19_in1_ready;

	assign branchC_19_clk = clk;
	assign branchC_19_rst = rst;
	assign Buffer_105_in1_data = branchC_19_out1_data;
	assign Buffer_105_in1_valid = branchC_19_out1_valid;
	assign branchC_19_out1_ready = Buffer_105_in1_ready;
	assign phiC_9_in1_data = branchC_19_out2_data;
	assign phiC_9_in1_valid = branchC_19_out2_valid;
	assign branchC_19_out2_ready = phiC_9_in1_ready;

	assign fork_28_clk = clk;
	assign fork_28_rst = rst;
	assign branch_7_in2_data = fork_28_out1_data;
	assign branch_7_in2_valid = fork_28_out1_valid;
	assign fork_28_out1_ready = branch_7_in2_ready;
	assign branchC_19_in2_data = fork_28_out2_data;
	assign branchC_19_in2_valid = fork_28_out2_valid;
	assign fork_28_out2_ready = branchC_19_in2_ready;

	assign source_3_clk = clk;
	assign source_3_rst = rst;
	assign cst_5_in1_data = source_3_out1_data;
	assign cst_5_in1_valid = source_3_out1_valid;
	assign source_3_out1_ready = cst_5_in1_ready;

	assign source_4_clk = clk;
	assign source_4_rst = rst;
	assign cst_6_in1_data = source_4_out1_data;
	assign cst_6_in1_valid = source_4_out1_valid;
	assign source_4_out1_ready = cst_6_in1_ready;

	assign ret_0_clk = clk;
	assign ret_0_rst = rst;
	assign end_0_in6_data = ret_0_out1_data;
	assign end_0_in6_valid = ret_0_out1_valid;
	assign ret_0_out1_ready = end_0_in6_ready;

	assign end_0_clk = clk;
	assign end_0_rst = rst;
	assign end_out = end_0_out1_data;
	assign end_0_out1_ready = end_ready;
	assign end_valid = end_0_out1_valid;

	assign phiC_13_clk = clk;
	assign phiC_13_rst = rst;
	assign ret_0_in1_data = phiC_13_out1_data;
	assign ret_0_in1_valid = phiC_13_out1_valid;
	assign phiC_13_out1_ready = ret_0_in1_ready;

	assign MC_x1_clk = clk;
	assign MC_x1_rst = rst;
	assign x1_ce0 = x1_we0;
	assign load_4_in1_data = MC_x1_out1_data;
	assign load_4_in1_valid = MC_x1_out1_valid;
	assign MC_x1_out1_ready = load_4_in1_ready;
	assign end_0_in1_data = MC_x1_out2_data;
	assign end_0_in1_valid = MC_x1_out2_valid;
	assign MC_x1_out2_ready = end_0_in1_ready;

	assign MC_A_clk = clk;
	assign MC_A_rst = rst;
	assign A_ce0 = A_we0;
	assign MC_A_in3_valid = 0;
	assign MC_A_in3_data = 0;
	assign load_12_in1_data = MC_A_out1_data;
	assign load_12_in1_valid = MC_A_out1_valid;
	assign MC_A_out1_ready = load_12_in1_ready;
	assign load_38_in1_data = MC_A_out2_data;
	assign load_38_in1_valid = MC_A_out2_valid;
	assign MC_A_out2_ready = load_38_in1_ready;
	assign end_0_in2_data = MC_A_out3_data;
	assign end_0_in2_valid = MC_A_out3_valid;
	assign MC_A_out3_ready = end_0_in2_ready;

	assign MC_y1_clk = clk;
	assign MC_y1_rst = rst;
	assign y1_ce0 = y1_we0;
	assign MC_y1_in2_valid = 0;
	assign MC_y1_in2_data = 0;
	assign load_15_in1_data = MC_y1_out1_data;
	assign load_15_in1_valid = MC_y1_out1_valid;
	assign MC_y1_out1_ready = load_15_in1_ready;
	assign end_0_in3_data = MC_y1_out2_data;
	assign end_0_in3_valid = MC_y1_out2_valid;
	assign MC_y1_out2_ready = end_0_in3_ready;

	assign MC_x2_clk = clk;
	assign MC_x2_rst = rst;
	assign x2_ce0 = x2_we0;
	assign load_30_in1_data = MC_x2_out1_data;
	assign load_30_in1_valid = MC_x2_out1_valid;
	assign MC_x2_out1_ready = load_30_in1_ready;
	assign end_0_in4_data = MC_x2_out2_data;
	assign end_0_in4_valid = MC_x2_out2_valid;
	assign MC_x2_out2_ready = end_0_in4_ready;

	assign MC_y2_clk = clk;
	assign MC_y2_rst = rst;
	assign y2_ce0 = y2_we0;
	assign MC_y2_in2_valid = 0;
	assign MC_y2_in2_data = 0;
	assign load_41_in1_data = MC_y2_out1_data;
	assign load_41_in1_valid = MC_y2_out1_valid;
	assign MC_y2_out1_ready = load_41_in1_ready;
	assign end_0_in5_data = MC_y2_out2_data;
	assign end_0_in5_valid = MC_y2_out2_valid;
	assign MC_y2_out2_ready = end_0_in5_ready;

	assign sink_0_clk = clk;
	assign sink_0_rst = rst;

	assign sink_1_clk = clk;
	assign sink_1_rst = rst;

	assign sink_2_clk = clk;
	assign sink_2_rst = rst;

	assign sink_3_clk = clk;
	assign sink_3_rst = rst;

	assign sink_4_clk = clk;
	assign sink_4_rst = rst;

	assign sink_5_clk = clk;
	assign sink_5_rst = rst;

	assign sink_6_clk = clk;
	assign sink_6_rst = rst;

	assign sink_7_clk = clk;
	assign sink_7_rst = rst;

	assign sink_8_clk = clk;
	assign sink_8_rst = rst;

	assign sink_9_clk = clk;
	assign sink_9_rst = rst;

	assign sink_10_clk = clk;
	assign sink_10_rst = rst;

	assign sink_11_clk = clk;
	assign sink_11_rst = rst;

	assign sink_12_clk = clk;
	assign sink_12_rst = rst;

	assign sink_13_clk = clk;
	assign sink_13_rst = rst;

	assign sink_14_clk = clk;
	assign sink_14_rst = rst;

	assign sink_15_clk = clk;
	assign sink_15_rst = rst;

	assign Buffer_100_clk = clk;
	assign Buffer_100_rst = rst;
	assign phi_6_in3_data = Buffer_100_out1_data;
	assign phi_6_in3_valid = Buffer_100_out1_valid;
	assign Buffer_100_out1_ready = phi_6_in3_ready;

	assign Buffer_101_clk = clk;
	assign Buffer_101_rst = rst;
	assign phi_7_in3_data = Buffer_101_out1_data;
	assign phi_7_in3_valid = Buffer_101_out1_valid;
	assign Buffer_101_out1_ready = phi_7_in3_ready;

	assign Buffer_102_clk = clk;
	assign Buffer_102_rst = rst;
	assign phi_n2_in2_data = Buffer_102_out1_data;
	assign phi_n2_in2_valid = Buffer_102_out1_valid;
	assign Buffer_102_out1_ready = phi_n2_in2_ready;

	assign Buffer_103_clk = clk;
	assign Buffer_103_rst = rst;
	assign phiC_7_in2_data = Buffer_103_out1_data;
	assign phiC_7_in2_valid = Buffer_103_out1_valid;
	assign Buffer_103_out1_ready = phiC_7_in2_ready;

	assign Buffer_104_clk = clk;
	assign Buffer_104_rst = rst;
	assign phi_1_in3_data = Buffer_104_out1_data;
	assign phi_1_in3_valid = Buffer_104_out1_valid;
	assign Buffer_104_out1_ready = phi_1_in3_ready;

	assign Buffer_105_clk = clk;
	assign Buffer_105_rst = rst;
	assign phiC_6_in2_data = Buffer_105_out1_data;
	assign phiC_6_in2_valid = Buffer_105_out1_valid;
	assign Buffer_105_out1_ready = phiC_6_in2_ready;

	assign Buffer_106_clk = clk;
	assign Buffer_106_rst = rst;
	assign phi_32_in3_data = Buffer_106_out1_data;
	assign phi_32_in3_valid = Buffer_106_out1_valid;
	assign Buffer_106_out1_ready = phi_32_in3_ready;

	assign Buffer_107_clk = clk;
	assign Buffer_107_rst = rst;
	assign phi_33_in3_data = Buffer_107_out1_data;
	assign phi_33_in3_valid = Buffer_107_out1_valid;
	assign Buffer_107_out1_ready = phi_33_in3_ready;

	assign Buffer_108_clk = clk;
	assign Buffer_108_rst = rst;
	assign phi_n5_in2_data = Buffer_108_out1_data;
	assign phi_n5_in2_valid = Buffer_108_out1_valid;
	assign Buffer_108_out1_ready = phi_n5_in2_ready;

	assign Buffer_109_clk = clk;
	assign Buffer_109_rst = rst;
	assign phiC_11_in2_data = Buffer_109_out1_data;
	assign phiC_11_in2_valid = Buffer_109_out1_valid;
	assign Buffer_109_out1_ready = phiC_11_in2_ready;

	assign Buffer_110_clk = clk;
	assign Buffer_110_rst = rst;
	assign phi_27_in3_data = Buffer_110_out1_data;
	assign phi_27_in3_valid = Buffer_110_out1_valid;
	assign Buffer_110_out1_ready = phi_27_in3_ready;

	assign Buffer_111_clk = clk;
	assign Buffer_111_rst = rst;
	assign phiC_10_in2_data = Buffer_111_out1_data;
	assign phiC_10_in2_valid = Buffer_111_out1_valid;
	assign Buffer_111_out1_ready = phiC_10_in2_ready;

	assign and_300_clk = clk;
	assign and_300_rst = rst;
	assign Buffer_300_in1_data = and_300_out1_data;
	assign Buffer_300_in1_valid = and_300_out1_valid;
	assign and_300_out1_ready = Buffer_300_in1_ready;

	assign Buffer_300_clk = clk;
	assign Buffer_300_rst = rst;
	assign and_301_in2_data = Buffer_300_out1_data;
	assign and_301_in2_valid = Buffer_300_out1_valid;
	assign Buffer_300_out1_ready = and_301_in2_ready;

	assign and_301_clk = clk;
	assign and_301_rst = rst;
	assign Buffer_301_in1_data = and_301_out1_data;
	assign Buffer_301_in1_valid = and_301_out1_valid;
	assign and_301_out1_ready = Buffer_301_in1_ready;

	assign Buffer_301_clk = clk;
	assign Buffer_301_rst = rst;
	assign branch_4_in1_data = Buffer_301_out1_data;
	assign branch_4_in1_valid = Buffer_301_out1_valid;
	assign Buffer_301_out1_ready = branch_4_in1_ready;

	assign and_302_clk = clk;
	assign and_302_rst = rst;
	assign Buffer_302_in1_data = and_302_out1_data;
	assign Buffer_302_in1_valid = and_302_out1_valid;
	assign and_302_out1_ready = Buffer_302_in1_ready;

	assign Buffer_302_clk = clk;
	assign Buffer_302_rst = rst;
	assign and_303_in2_data = Buffer_302_out1_data;
	assign and_303_in2_valid = Buffer_302_out1_valid;
	assign Buffer_302_out1_ready = and_303_in2_ready;

	assign and_303_clk = clk;
	assign and_303_rst = rst;
	assign Buffer_303_in1_data = and_303_out1_data;
	assign Buffer_303_in1_valid = and_303_out1_valid;
	assign and_303_out1_ready = Buffer_303_in1_ready;

	assign Buffer_303_clk = clk;
	assign Buffer_303_rst = rst;
	assign branch_12_in1_data = Buffer_303_out1_data;
	assign branch_12_in1_valid = Buffer_303_out1_valid;
	assign Buffer_303_out1_ready = branch_12_in1_ready;

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_1
		(.clk(phi_1_clk), .rst(phi_1_rst),
		.data_in_bus({{5'b0, phi_1_in1_data}, phi_1_in3_data, phi_1_in2_data}), .valid_in_bus({phi_1_in1_valid, phi_1_in3_valid, phi_1_in2_valid}), .ready_in_bus({phi_1_in1_ready, phi_1_in3_ready, phi_1_in2_ready}), 
		.data_out_bus({phi_1_out1_data}), .valid_out_bus({phi_1_out1_valid}), .ready_out_bus({phi_1_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_4
		(.clk(load_4_clk), .rst(load_4_rst),
		.data_in_bus({load_4_in1_data}), .address_in_bus({load_4_in2_data}), .valid_in_bus({load_4_in2_valid, load_4_in1_valid}), .ready_in_bus({load_4_in2_ready, load_4_in1_ready}), 
		.data_out_bus({load_4_out1_data}), .address_out_bus({load_4_out2_data}), .valid_out_bus({load_4_out2_valid, load_4_out1_valid}), .ready_out_bus({load_4_out2_ready, load_4_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block2
		(.clk(brCst_block2_clk), .rst(brCst_block2_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block2_in1_valid}), .ready_in_bus({brCst_block2_in1_ready}), 
		.data_out_bus({brCst_block2_out1_data}), .valid_out_bus({brCst_block2_out1_valid}), .ready_out_bus({brCst_block2_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_1
		(.clk(cst_1_clk), .rst(cst_1_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_1_in1_valid}), .ready_in_bus({cst_1_in1_ready}), 
		.data_out_bus({cst_1_out1_data}), .valid_out_bus({cst_1_out1_valid}), .ready_out_bus({cst_1_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_0
		(.clk(fork_0_clk), .rst(fork_0_rst),
		.data_in_bus({fork_0_in1_data}), .valid_in_bus({fork_0_in1_valid}), .ready_in_bus({fork_0_in1_ready}), 
		.data_out_bus({fork_0_out2_data, fork_0_out1_data}), .valid_out_bus({fork_0_out2_valid, fork_0_out1_valid}), .ready_out_bus({fork_0_out2_ready, fork_0_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_1
		(.clk(branch_1_clk), .rst(branch_1_rst),
		.data_in_bus({{31'b0, branch_1_in2_data}, branch_1_in1_data}), .valid_in_bus({branch_1_in2_valid, branch_1_in1_valid}), .ready_in_bus({branch_1_in2_ready, branch_1_in1_ready}), 
		.data_out_bus({branch_1_out2_data, branch_1_out1_data}), .valid_out_bus({branch_1_out2_valid, branch_1_out1_valid}), .ready_out_bus({branch_1_out2_ready, branch_1_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_2
		(.clk(branch_2_clk), .rst(branch_2_rst),
		.data_in_bus({{branch_2_in2_data}, branch_2_in1_data}), .valid_in_bus({branch_2_in2_valid, branch_2_in1_valid}), .ready_in_bus({branch_2_in2_ready, branch_2_in1_ready}), 
		.data_out_bus({branch_2_out2_data, branch_2_out1_data}), .valid_out_bus({branch_2_out2_valid, branch_2_out1_valid}), .ready_out_bus({branch_2_out2_ready, branch_2_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_3
		(.clk(branch_3_clk), .rst(branch_3_rst),
		.data_in_bus({{5'b0, branch_3_in2_data}, branch_3_in1_data}), .valid_in_bus({branch_3_in2_valid, branch_3_in1_valid}), .ready_in_bus({branch_3_in2_ready, branch_3_in1_ready}), 
		.data_out_bus({branch_3_out2_data, branch_3_out1_data}), .valid_out_bus({branch_3_out2_valid, branch_3_out1_valid}), .ready_out_bus({branch_3_out2_ready, branch_3_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_15
		(.clk(fork_15_clk), .rst(fork_15_rst),
		.data_in_bus({fork_15_in1_data}), .valid_in_bus({fork_15_in1_valid}), .ready_in_bus({fork_15_in1_ready}), 
		.data_out_bus({fork_15_out4_data, fork_15_out3_data, fork_15_out2_data, fork_15_out1_data}), .valid_out_bus({fork_15_out4_valid, fork_15_out3_valid, fork_15_out2_valid, fork_15_out1_valid}), .ready_out_bus({fork_15_out4_ready, fork_15_out3_ready, fork_15_out2_ready, fork_15_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_6
		(.clk(phiC_6_clk), .rst(phiC_6_rst),
		.data_in_bus({phiC_6_in2_data, phiC_6_in1_data}), .valid_in_bus({phiC_6_in2_valid, phiC_6_in1_valid}), .ready_in_bus({phiC_6_in2_ready, phiC_6_in1_ready}), 
		.data_out_bus({phiC_6_out2_data, phiC_6_out1_data}), .valid_out_bus({phiC_6_out2_valid, phiC_6_out1_valid}), .ready_out_bus({phiC_6_out2_ready, phiC_6_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_25
		(.clk(forkC_25_clk), .rst(forkC_25_rst),
		.data_in_bus({forkC_25_in1_data}), .valid_in_bus({forkC_25_in1_valid}), .ready_in_bus({forkC_25_in1_ready}), 
		.data_out_bus({forkC_25_out3_data, forkC_25_out2_data, forkC_25_out1_data}), .valid_out_bus({forkC_25_out3_valid, forkC_25_out2_valid, forkC_25_out1_valid}), .ready_out_bus({forkC_25_out3_ready, forkC_25_out2_ready, forkC_25_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_17
		(.clk(branchC_17_clk), .rst(branchC_17_rst),
		.data_in_bus({{branchC_17_in2_data}, branchC_17_in1_data}), .valid_in_bus({branchC_17_in2_valid, branchC_17_in1_valid}), .ready_in_bus({branchC_17_in2_ready, branchC_17_in1_ready}), 
		.data_out_bus({branchC_17_out2_data, branchC_17_out1_data}), .valid_out_bus({branchC_17_out2_valid, branchC_17_out1_valid}), .ready_out_bus({branchC_17_out2_ready, branchC_17_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block1
		(.clk(brCst_block1_clk), .rst(brCst_block1_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block1_in1_valid}), .ready_in_bus({brCst_block1_in1_ready}), 
		.data_out_bus({brCst_block1_out1_data}), .valid_out_bus({brCst_block1_out1_valid}), .ready_out_bus({brCst_block1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_0
		(.clk(cst_0_clk), .rst(cst_0_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_0_in1_valid}), .ready_in_bus({cst_0_in1_ready}), 
		.data_out_bus({cst_0_out1_data}), .valid_out_bus({cst_0_out1_valid}), .ready_out_bus({cst_0_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_0
		(.clk(branch_0_clk), .rst(branch_0_rst),
		.data_in_bus({{branch_0_in2_data}, branch_0_in1_data}), .valid_in_bus({branch_0_in2_valid, branch_0_in1_valid}), .ready_in_bus({branch_0_in2_ready, branch_0_in1_ready}), 
		.data_out_bus({branch_0_out2_data, branch_0_out1_data}), .valid_out_bus({branch_0_out2_valid, branch_0_out1_valid}), .ready_out_bus({branch_0_out2_ready, branch_0_out1_ready}));

	start_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) start_node_start_0
		(.clk(start_0_clk), .rst(start_0_rst),
		.data_in_bus({start_0_in1_data}), .valid_in_bus({start_0_in1_valid}), .ready_in_bus({start_0_in1_ready}), 
		.data_out_bus({start_0_out1_data}), .valid_out_bus({start_0_out1_valid}), .ready_out_bus({start_0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_23
		(.clk(forkC_23_clk), .rst(forkC_23_rst),
		.data_in_bus({forkC_23_in1_data}), .valid_in_bus({forkC_23_in1_valid}), .ready_in_bus({forkC_23_in1_ready}), 
		.data_out_bus({forkC_23_out3_data, forkC_23_out2_data, forkC_23_out1_data}), .valid_out_bus({forkC_23_out3_valid, forkC_23_out2_valid, forkC_23_out1_valid}), .ready_out_bus({forkC_23_out3_ready, forkC_23_out2_ready, forkC_23_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_16
		(.clk(branchC_16_clk), .rst(branchC_16_rst),
		.data_in_bus({{branchC_16_in2_data}, branchC_16_in1_data}), .valid_in_bus({branchC_16_in2_valid, branchC_16_in1_valid}), .ready_in_bus({branchC_16_in2_ready, branchC_16_in1_ready}), 
		.data_out_bus({branchC_16_out2_data, branchC_16_out1_data}), .valid_out_bus({branchC_16_out2_valid, branchC_16_out1_valid}), .ready_out_bus({branchC_16_out2_ready, branchC_16_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_24
		(.clk(fork_24_clk), .rst(fork_24_rst),
		.data_in_bus({fork_24_in1_data}), .valid_in_bus({fork_24_in1_valid}), .ready_in_bus({fork_24_in1_ready}), 
		.data_out_bus({fork_24_out2_data, fork_24_out1_data}), .valid_out_bus({fork_24_out2_valid, fork_24_out1_valid}), .ready_out_bus({fork_24_out2_ready, fork_24_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_27
		(.clk(phi_27_clk), .rst(phi_27_rst),
		.data_in_bus({{5'b0, phi_27_in1_data}, phi_27_in3_data, phi_27_in2_data}), .valid_in_bus({phi_27_in1_valid, phi_27_in3_valid, phi_27_in2_valid}), .ready_in_bus({phi_27_in1_ready, phi_27_in3_ready, phi_27_in2_ready}), 
		.data_out_bus({phi_27_out1_data}), .valid_out_bus({phi_27_out1_valid}), .ready_out_bus({phi_27_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_30
		(.clk(load_30_clk), .rst(load_30_rst),
		.data_in_bus({load_30_in1_data}), .address_in_bus({load_30_in2_data}), .valid_in_bus({load_30_in2_valid, load_30_in1_valid}), .ready_in_bus({load_30_in2_ready, load_30_in1_ready}), 
		.data_out_bus({load_30_out1_data}), .address_out_bus({load_30_out2_data}), .valid_out_bus({load_30_out2_valid, load_30_out1_valid}), .ready_out_bus({load_30_out2_ready, load_30_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block6
		(.clk(brCst_block6_clk), .rst(brCst_block6_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block6_in1_valid}), .ready_in_bus({brCst_block6_in1_ready}), 
		.data_out_bus({brCst_block6_out1_data}), .valid_out_bus({brCst_block6_out1_valid}), .ready_out_bus({brCst_block6_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_8
		(.clk(cst_8_clk), .rst(cst_8_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_8_in1_valid}), .ready_in_bus({cst_8_in1_ready}), 
		.data_out_bus({cst_8_out1_data}), .valid_out_bus({cst_8_out1_valid}), .ready_out_bus({cst_8_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_5
		(.clk(fork_5_clk), .rst(fork_5_rst),
		.data_in_bus({fork_5_in1_data}), .valid_in_bus({fork_5_in1_valid}), .ready_in_bus({fork_5_in1_ready}), 
		.data_out_bus({fork_5_out2_data, fork_5_out1_data}), .valid_out_bus({fork_5_out2_valid, fork_5_out1_valid}), .ready_out_bus({fork_5_out2_ready, fork_5_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_9
		(.clk(branch_9_clk), .rst(branch_9_rst),
		.data_in_bus({{31'b0, branch_9_in2_data}, branch_9_in1_data}), .valid_in_bus({branch_9_in2_valid, branch_9_in1_valid}), .ready_in_bus({branch_9_in2_ready, branch_9_in1_ready}), 
		.data_out_bus({branch_9_out2_data, branch_9_out1_data}), .valid_out_bus({branch_9_out2_valid, branch_9_out1_valid}), .ready_out_bus({branch_9_out2_ready, branch_9_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_10
		(.clk(branch_10_clk), .rst(branch_10_rst),
		.data_in_bus({{branch_10_in2_data}, branch_10_in1_data}), .valid_in_bus({branch_10_in2_valid, branch_10_in1_valid}), .ready_in_bus({branch_10_in2_ready, branch_10_in1_ready}), 
		.data_out_bus({branch_10_out2_data, branch_10_out1_data}), .valid_out_bus({branch_10_out2_valid, branch_10_out1_valid}), .ready_out_bus({branch_10_out2_ready, branch_10_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_11
		(.clk(branch_11_clk), .rst(branch_11_rst),
		.data_in_bus({{5'b0, branch_11_in2_data}, branch_11_in1_data}), .valid_in_bus({branch_11_in2_valid, branch_11_in1_valid}), .ready_in_bus({branch_11_in2_ready, branch_11_in1_ready}), 
		.data_out_bus({branch_11_out2_data, branch_11_out1_data}), .valid_out_bus({branch_11_out2_valid, branch_11_out1_valid}), .ready_out_bus({branch_11_out2_ready, branch_11_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_19
		(.clk(fork_19_clk), .rst(fork_19_rst),
		.data_in_bus({fork_19_in1_data}), .valid_in_bus({fork_19_in1_valid}), .ready_in_bus({fork_19_in1_ready}), 
		.data_out_bus({fork_19_out4_data, fork_19_out3_data, fork_19_out2_data, fork_19_out1_data}), .valid_out_bus({fork_19_out4_valid, fork_19_out3_valid, fork_19_out2_valid, fork_19_out1_valid}), .ready_out_bus({fork_19_out4_ready, fork_19_out3_ready, fork_19_out2_ready, fork_19_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_10
		(.clk(phiC_10_clk), .rst(phiC_10_rst),
		.data_in_bus({phiC_10_in2_data, phiC_10_in1_data}), .valid_in_bus({phiC_10_in2_valid, phiC_10_in1_valid}), .ready_in_bus({phiC_10_in2_ready, phiC_10_in1_ready}), 
		.data_out_bus({phiC_10_out2_data, phiC_10_out1_data}), .valid_out_bus({phiC_10_out2_valid, phiC_10_out1_valid}), .ready_out_bus({phiC_10_out2_ready, phiC_10_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_31
		(.clk(forkC_31_clk), .rst(forkC_31_rst),
		.data_in_bus({forkC_31_in1_data}), .valid_in_bus({forkC_31_in1_valid}), .ready_in_bus({forkC_31_in1_ready}), 
		.data_out_bus({forkC_31_out3_data, forkC_31_out2_data, forkC_31_out1_data}), .valid_out_bus({forkC_31_out3_valid, forkC_31_out2_valid, forkC_31_out1_valid}), .ready_out_bus({forkC_31_out3_ready, forkC_31_out2_ready, forkC_31_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_21
		(.clk(branchC_21_clk), .rst(branchC_21_rst),
		.data_in_bus({{branchC_21_in2_data}, branchC_21_in1_data}), .valid_in_bus({branchC_21_in2_valid, branchC_21_in1_valid}), .ready_in_bus({branchC_21_in2_ready, branchC_21_in1_ready}), 
		.data_out_bus({branchC_21_out2_data, branchC_21_out1_data}), .valid_out_bus({branchC_21_out2_valid, branchC_21_out1_valid}), .ready_out_bus({branchC_21_out2_ready, branchC_21_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_32
		(.clk(phi_32_clk), .rst(phi_32_rst),
		.data_in_bus({{31'b0, phi_32_in1_data}, phi_32_in3_data, phi_32_in2_data}), .valid_in_bus({phi_32_in1_valid, phi_32_in3_valid, phi_32_in2_valid}), .ready_in_bus({phi_32_in1_ready, phi_32_in3_ready, phi_32_in2_ready}), 
		.data_out_bus({phi_32_out1_data}), .valid_out_bus({phi_32_out1_valid}), .ready_out_bus({phi_32_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_33
		(.clk(phi_33_clk), .rst(phi_33_rst),
		.data_in_bus({{5'b0, phi_33_in1_data}, phi_33_in3_data, phi_33_in2_data}), .valid_in_bus({phi_33_in1_valid, phi_33_in3_valid, phi_33_in2_valid}), .ready_in_bus({phi_33_in1_ready, phi_33_in3_ready, phi_33_in2_ready}), 
		.data_out_bus({phi_33_out1_data}), .valid_out_bus({phi_33_out1_valid}), .ready_out_bus({phi_33_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_9
		(.clk(cst_9_clk), .rst(cst_9_rst),
		.data_in_bus({3'd5}), .valid_in_bus({cst_9_in1_valid}), .ready_in_bus({cst_9_in1_ready}), 
		.data_out_bus({cst_9_out1_data}), .valid_out_bus({cst_9_out1_valid}), .ready_out_bus({cst_9_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(11), .DATA_OUT_SIZE(11)) shl_op_shl_34
		(.clk(shl_34_clk), .rst(shl_34_rst),
		.data_in_bus({shl_34_in2_data, shl_34_in1_data}), .valid_in_bus({shl_34_in2_valid, shl_34_in1_valid}), .ready_in_bus({shl_34_in2_ready, shl_34_in1_ready}), 
		.data_out_bus({shl_34_out1_data}), .valid_out_bus({shl_34_out1_valid}), .ready_out_bus({shl_34_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(12), .DATA_OUT_SIZE(12)) add_op_add_35
		(.clk(add_35_clk), .rst(add_35_rst),
		.data_in_bus({add_35_in2_data, add_35_in1_data}), .valid_in_bus({add_35_in2_valid, add_35_in1_valid}), .ready_in_bus({add_35_in2_ready, add_35_in1_ready}), 
		.data_out_bus({add_35_out1_data}), .valid_out_bus({add_35_out1_valid}), .ready_out_bus({add_35_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(12), .DATA_SIZE(32)) mc_load_op_load_38
		(.clk(load_38_clk), .rst(load_38_rst),
		.data_in_bus({load_38_in1_data}), .address_in_bus({load_38_in2_data}), .valid_in_bus({load_38_in2_valid, load_38_in1_valid}), .ready_in_bus({load_38_in2_ready, load_38_in1_ready}), 
		.data_out_bus({load_38_out1_data}), .address_out_bus({load_38_out2_data}), .valid_out_bus({load_38_out2_valid, load_38_out1_valid}), .ready_out_bus({load_38_out2_ready, load_38_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_41
		(.clk(load_41_clk), .rst(load_41_rst),
		.data_in_bus({load_41_in1_data}), .address_in_bus({load_41_in2_data}), .valid_in_bus({load_41_in2_valid, load_41_in1_valid}), .ready_in_bus({load_41_in2_ready, load_41_in1_ready}), 
		.data_out_bus({load_41_out1_data}), .address_out_bus({load_41_out2_data}), .valid_out_bus({load_41_out2_valid, load_41_out1_valid}), .ready_out_bus({load_41_out2_ready, load_41_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_10
		(.clk(cst_10_clk), .rst(cst_10_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_10_in1_valid}), .ready_in_bus({cst_10_in1_ready}), 
		.data_out_bus({cst_10_out1_data}), .valid_out_bus({cst_10_out1_valid}), .ready_out_bus({cst_10_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_44
		(.clk(add_44_clk), .rst(add_44_rst),
		.data_in_bus({add_44_in2_data, add_44_in1_data}), .valid_in_bus({add_44_in2_valid, add_44_in1_valid}), .ready_in_bus({add_44_in2_ready, add_44_in1_ready}), 
		.data_out_bus({add_44_out1_data}), .valid_out_bus({add_44_out1_valid}), .ready_out_bus({add_44_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_11
		(.clk(cst_11_clk), .rst(cst_11_rst),
		.data_in_bus({6'd32}), .valid_in_bus({cst_11_in1_valid}), .ready_in_bus({cst_11_in1_ready}), 
		.data_out_bus({cst_11_out1_data}), .valid_out_bus({cst_11_out1_valid}), .ready_out_bus({cst_11_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_45
		(.clk(icmp_45_clk), .rst(icmp_45_rst),
		.data_in_bus({icmp_45_in2_data, icmp_45_in1_data}), .valid_in_bus({icmp_45_in2_valid, icmp_45_in1_valid}), .ready_in_bus({icmp_45_in2_ready, icmp_45_in1_ready}), 
		.data_out_bus({icmp_45_out1_data}), .valid_out_bus({icmp_45_out1_valid}), .ready_out_bus({icmp_45_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n5
		(.clk(phi_n5_clk), .rst(phi_n5_rst),
		.data_in_bus({phi_n5_in2_data, phi_n5_in1_data}), .valid_in_bus({phi_n5_in2_valid, phi_n5_in1_valid}), .ready_in_bus({phi_n5_in2_ready, phi_n5_in1_ready}), 
		.data_out_bus({phi_n5_out1_data}), .valid_out_bus({phi_n5_out1_valid}), .ready_out_bus({phi_n5_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_6
		(.clk(fork_6_clk), .rst(fork_6_rst),
		.data_in_bus({fork_6_in1_data}), .valid_in_bus({fork_6_in1_valid}), .ready_in_bus({fork_6_in1_ready}), 
		.data_out_bus({fork_6_out3_data, fork_6_out2_data, fork_6_out1_data}), .valid_out_bus({fork_6_out3_valid, fork_6_out2_valid, fork_6_out1_valid}), .ready_out_bus({fork_6_out3_ready, fork_6_out2_ready, fork_6_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_8
		(.clk(fork_8_clk), .rst(fork_8_rst),
		.data_in_bus({fork_8_in1_data}), .valid_in_bus({fork_8_in1_valid}), .ready_in_bus({fork_8_in1_ready}), 
		.data_out_bus({fork_8_out2_data, fork_8_out1_data}), .valid_out_bus({fork_8_out2_valid, fork_8_out1_valid}), .ready_out_bus({fork_8_out2_ready, fork_8_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_13
		(.clk(fork_13_clk), .rst(fork_13_rst),
		.data_in_bus({fork_13_in1_data}), .valid_in_bus({fork_13_in1_valid}), .ready_in_bus({fork_13_in1_ready}), 
		.data_out_bus({fork_13_out2_data, fork_13_out1_data}), .valid_out_bus({fork_13_out2_valid, fork_13_out1_valid}), .ready_out_bus({fork_13_out2_ready, fork_13_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_12
		(.clk(branch_12_clk), .rst(branch_12_rst),
		.data_in_bus({{31'b0, branch_12_in2_data}, branch_12_in1_data}), .valid_in_bus({branch_12_in2_valid, branch_12_in1_valid}), .ready_in_bus({branch_12_in2_ready, branch_12_in1_ready}), 
		.data_out_bus({branch_12_out2_data, branch_12_out1_data}), .valid_out_bus({branch_12_out2_valid, branch_12_out1_valid}), .ready_out_bus({branch_12_out2_ready, branch_12_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_13
		(.clk(branch_13_clk), .rst(branch_13_rst),
		.data_in_bus({{5'b0, branch_13_in2_data}, branch_13_in1_data}), .valid_in_bus({branch_13_in2_valid, branch_13_in1_valid}), .ready_in_bus({branch_13_in2_ready, branch_13_in1_ready}), 
		.data_out_bus({branch_13_out2_data, branch_13_out1_data}), .valid_out_bus({branch_13_out2_valid, branch_13_out1_valid}), .ready_out_bus({branch_13_out2_ready, branch_13_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_14
		(.clk(branch_14_clk), .rst(branch_14_rst),
		.data_in_bus({{5'b0, branch_14_in2_data}, branch_14_in1_data}), .valid_in_bus({branch_14_in2_valid, branch_14_in1_valid}), .ready_in_bus({branch_14_in2_ready, branch_14_in1_ready}), 
		.data_out_bus({branch_14_out2_data, branch_14_out1_data}), .valid_out_bus({branch_14_out2_valid, branch_14_out1_valid}), .ready_out_bus({branch_14_out2_ready, branch_14_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_20
		(.clk(fork_20_clk), .rst(fork_20_rst),
		.data_in_bus({fork_20_in1_data}), .valid_in_bus({fork_20_in1_valid}), .ready_in_bus({fork_20_in1_ready}), 
		.data_out_bus({fork_20_out4_data, fork_20_out3_data, fork_20_out2_data, fork_20_out1_data}), .valid_out_bus({fork_20_out4_valid, fork_20_out3_valid, fork_20_out2_valid, fork_20_out1_valid}), .ready_out_bus({fork_20_out4_ready, fork_20_out3_ready, fork_20_out2_ready, fork_20_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_11
		(.clk(phiC_11_clk), .rst(phiC_11_rst),
		.data_in_bus({phiC_11_in2_data, phiC_11_in1_data}), .valid_in_bus({phiC_11_in2_valid, phiC_11_in1_valid}), .ready_in_bus({phiC_11_in2_ready, phiC_11_in1_ready}), 
		.data_out_bus({phiC_11_out2_data, phiC_11_out1_data}), .valid_out_bus({phiC_11_out2_valid, phiC_11_out1_valid}), .ready_out_bus({phiC_11_out2_ready, phiC_11_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_22
		(.clk(branchC_22_clk), .rst(branchC_22_rst),
		.data_in_bus({{branchC_22_in2_data}, branchC_22_in1_data}), .valid_in_bus({branchC_22_in2_valid, branchC_22_in1_valid}), .ready_in_bus({branchC_22_in2_ready, branchC_22_in1_ready}), 
		.data_out_bus({branchC_22_out2_data, branchC_22_out1_data}), .valid_out_bus({branchC_22_out2_valid, branchC_22_out1_valid}), .ready_out_bus({branchC_22_out2_ready, branchC_22_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_5
		(.clk(source_5_clk), .rst(source_5_rst),
		.data_out_bus({source_5_out1_data}), .valid_out_bus({source_5_out1_valid}), .ready_out_bus({source_5_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_6
		(.clk(source_6_clk), .rst(source_6_rst),
		.data_out_bus({source_6_out1_data}), .valid_out_bus({source_6_out1_valid}), .ready_out_bus({source_6_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_7
		(.clk(source_7_clk), .rst(source_7_rst),
		.data_out_bus({source_7_out1_data}), .valid_out_bus({source_7_out1_valid}), .ready_out_bus({source_7_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_39
		(.clk(fork_39_clk), .rst(fork_39_rst),
		.data_in_bus({fork_39_in1_data}), .valid_in_bus({fork_39_in1_valid}), .ready_in_bus({fork_39_in1_ready}), 
		.data_out_bus({fork_39_out2_data, fork_39_out1_data}), .valid_out_bus({fork_39_out2_valid, fork_39_out1_valid}), .ready_out_bus({fork_39_out2_ready, fork_39_out1_ready}));

	mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_store_op_store_1
		(.clk(store_1_clk), .rst(store_1_rst),
		.data_in_bus({store_1_in1_data}), .address_in_bus({store_1_in2_data}), .valid_in_bus({store_1_in2_valid, store_1_in1_valid}), .ready_in_bus({store_1_in2_ready, store_1_in1_ready}), 
		.data_out_bus({store_1_out1_data}), .address_out_bus({store_1_out2_data}), .valid_out_bus({store_1_out2_valid, store_1_out1_valid}), .ready_out_bus({store_1_out2_ready, store_1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_12
		(.clk(cst_12_clk), .rst(cst_12_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_12_in1_valid}), .ready_in_bus({cst_12_in1_ready}), 
		.data_out_bus({cst_12_out1_data}), .valid_out_bus({cst_12_out1_valid}), .ready_out_bus({cst_12_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_49
		(.clk(add_49_clk), .rst(add_49_rst),
		.data_in_bus({add_49_in2_data, add_49_in1_data}), .valid_in_bus({add_49_in2_valid, add_49_in1_valid}), .ready_in_bus({add_49_in2_ready, add_49_in1_ready}), 
		.data_out_bus({add_49_out1_data}), .valid_out_bus({add_49_out1_valid}), .ready_out_bus({add_49_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_13
		(.clk(cst_13_clk), .rst(cst_13_rst),
		.data_in_bus({6'd32}), .valid_in_bus({cst_13_in1_valid}), .ready_in_bus({cst_13_in1_ready}), 
		.data_out_bus({cst_13_out1_data}), .valid_out_bus({cst_13_out1_valid}), .ready_out_bus({cst_13_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_50
		(.clk(icmp_50_clk), .rst(icmp_50_rst),
		.data_in_bus({icmp_50_in2_data, icmp_50_in1_data}), .valid_in_bus({icmp_50_in2_valid, icmp_50_in1_valid}), .ready_in_bus({icmp_50_in2_ready, icmp_50_in1_ready}), 
		.data_out_bus({icmp_50_out1_data}), .valid_out_bus({icmp_50_out1_valid}), .ready_out_bus({icmp_50_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n3
		(.clk(phi_n3_clk), .rst(phi_n3_rst),
		.data_in_bus({phi_n3_in1_data}), .valid_in_bus({phi_n3_in1_valid}), .ready_in_bus({phi_n3_in1_ready}), 
		.data_out_bus({phi_n3_out1_data}), .valid_out_bus({phi_n3_out1_valid}), .ready_out_bus({phi_n3_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n4
		(.clk(phi_n4_clk), .rst(phi_n4_rst),
		.data_in_bus({phi_n4_in1_data}), .valid_in_bus({phi_n4_in1_valid}), .ready_in_bus({phi_n4_in1_ready}), 
		.data_out_bus({phi_n4_out1_data}), .valid_out_bus({phi_n4_out1_valid}), .ready_out_bus({phi_n4_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_9
		(.clk(fork_9_clk), .rst(fork_9_rst),
		.data_in_bus({fork_9_in1_data}), .valid_in_bus({fork_9_in1_valid}), .ready_in_bus({fork_9_in1_ready}), 
		.data_out_bus({fork_9_out2_data, fork_9_out1_data}), .valid_out_bus({fork_9_out2_valid, fork_9_out1_valid}), .ready_out_bus({fork_9_out2_ready, fork_9_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_12
		(.clk(fork_12_clk), .rst(fork_12_rst),
		.data_in_bus({fork_12_in1_data}), .valid_in_bus({fork_12_in1_valid}), .ready_in_bus({fork_12_in1_ready}), 
		.data_out_bus({fork_12_out2_data, fork_12_out1_data}), .valid_out_bus({fork_12_out2_valid, fork_12_out1_valid}), .ready_out_bus({fork_12_out2_ready, fork_12_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_15
		(.clk(branch_15_clk), .rst(branch_15_rst),
		.data_in_bus({{5'b0, branch_15_in2_data}, branch_15_in1_data}), .valid_in_bus({branch_15_in2_valid, branch_15_in1_valid}), .ready_in_bus({branch_15_in2_ready, branch_15_in1_ready}), 
		.data_out_bus({branch_15_out2_data, branch_15_out1_data}), .valid_out_bus({branch_15_out2_valid, branch_15_out1_valid}), .ready_out_bus({branch_15_out2_ready, branch_15_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_15
		(.clk(cst_15_clk), .rst(cst_15_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_15_in1_valid}), .ready_in_bus({cst_15_in1_ready}), 
		.data_out_bus({cst_15_out1_data}), .valid_out_bus({cst_15_out1_valid}), .ready_out_bus({cst_15_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_12
		(.clk(phiC_12_clk), .rst(phiC_12_rst),
		.data_in_bus({phiC_12_in1_data}), .valid_in_bus({phiC_12_in1_valid}), .ready_in_bus({phiC_12_in1_ready}), 
		.data_out_bus({phiC_12_out1_data}), .valid_out_bus({phiC_12_out1_valid}), .ready_out_bus({phiC_12_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_33
		(.clk(forkC_33_clk), .rst(forkC_33_rst),
		.data_in_bus({forkC_33_in1_data}), .valid_in_bus({forkC_33_in1_valid}), .ready_in_bus({forkC_33_in1_ready}), 
		.data_out_bus({forkC_33_out2_data, forkC_33_out1_data}), .valid_out_bus({forkC_33_out2_valid, forkC_33_out1_valid}), .ready_out_bus({forkC_33_out2_ready, forkC_33_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_23
		(.clk(branchC_23_clk), .rst(branchC_23_rst),
		.data_in_bus({{branchC_23_in2_data}, branchC_23_in1_data}), .valid_in_bus({branchC_23_in2_valid, branchC_23_in1_valid}), .ready_in_bus({branchC_23_in2_ready, branchC_23_in1_ready}), 
		.data_out_bus({branchC_23_out2_data, branchC_23_out1_data}), .valid_out_bus({branchC_23_out2_valid, branchC_23_out1_valid}), .ready_out_bus({branchC_23_out2_ready, branchC_23_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_34
		(.clk(fork_34_clk), .rst(fork_34_rst),
		.data_in_bus({fork_34_in1_data}), .valid_in_bus({fork_34_in1_valid}), .ready_in_bus({fork_34_in1_ready}), 
		.data_out_bus({fork_34_out2_data, fork_34_out1_data}), .valid_out_bus({fork_34_out2_valid, fork_34_out1_valid}), .ready_out_bus({fork_34_out2_ready, fork_34_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_8
		(.clk(source_8_clk), .rst(source_8_rst),
		.data_out_bus({source_8_out1_data}), .valid_out_bus({source_8_out1_valid}), .ready_out_bus({source_8_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_9
		(.clk(source_9_clk), .rst(source_9_rst),
		.data_out_bus({source_9_out1_data}), .valid_out_bus({source_9_out1_valid}), .ready_out_bus({source_9_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block5
		(.clk(brCst_block5_clk), .rst(brCst_block5_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block5_in1_valid}), .ready_in_bus({brCst_block5_in1_ready}), 
		.data_out_bus({brCst_block5_out1_data}), .valid_out_bus({brCst_block5_out1_valid}), .ready_out_bus({brCst_block5_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_7
		(.clk(cst_7_clk), .rst(cst_7_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_7_in1_valid}), .ready_in_bus({cst_7_in1_ready}), 
		.data_out_bus({cst_7_out1_data}), .valid_out_bus({cst_7_out1_valid}), .ready_out_bus({cst_7_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_8
		(.clk(branch_8_clk), .rst(branch_8_rst),
		.data_in_bus({{branch_8_in2_data}, branch_8_in1_data}), .valid_in_bus({branch_8_in2_valid, branch_8_in1_valid}), .ready_in_bus({branch_8_in2_ready, branch_8_in1_ready}), 
		.data_out_bus({branch_8_out2_data, branch_8_out1_data}), .valid_out_bus({branch_8_out2_valid, branch_8_out1_valid}), .ready_out_bus({branch_8_out2_ready, branch_8_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_9
		(.clk(phiC_9_clk), .rst(phiC_9_rst),
		.data_in_bus({phiC_9_in1_data}), .valid_in_bus({phiC_9_in1_valid}), .ready_in_bus({phiC_9_in1_ready}), 
		.data_out_bus({phiC_9_out1_data}), .valid_out_bus({phiC_9_out1_valid}), .ready_out_bus({phiC_9_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_29
		(.clk(forkC_29_clk), .rst(forkC_29_rst),
		.data_in_bus({forkC_29_in1_data}), .valid_in_bus({forkC_29_in1_valid}), .ready_in_bus({forkC_29_in1_ready}), 
		.data_out_bus({forkC_29_out3_data, forkC_29_out2_data, forkC_29_out1_data}), .valid_out_bus({forkC_29_out3_valid, forkC_29_out2_valid, forkC_29_out1_valid}), .ready_out_bus({forkC_29_out3_ready, forkC_29_out2_ready, forkC_29_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_20
		(.clk(branchC_20_clk), .rst(branchC_20_rst),
		.data_in_bus({{branchC_20_in2_data}, branchC_20_in1_data}), .valid_in_bus({branchC_20_in2_valid, branchC_20_in1_valid}), .ready_in_bus({branchC_20_in2_ready, branchC_20_in1_ready}), 
		.data_out_bus({branchC_20_out2_data, branchC_20_out1_data}), .valid_out_bus({branchC_20_out2_valid, branchC_20_out1_valid}), .ready_out_bus({branchC_20_out2_ready, branchC_20_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_30
		(.clk(fork_30_clk), .rst(fork_30_rst),
		.data_in_bus({fork_30_in1_data}), .valid_in_bus({fork_30_in1_valid}), .ready_in_bus({fork_30_in1_ready}), 
		.data_out_bus({fork_30_out2_data, fork_30_out1_data}), .valid_out_bus({fork_30_out2_valid, fork_30_out1_valid}), .ready_out_bus({fork_30_out2_ready, fork_30_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_6
		(.clk(phi_6_clk), .rst(phi_6_rst),
		.data_in_bus({{31'b0, phi_6_in1_data}, phi_6_in3_data, phi_6_in2_data}), .valid_in_bus({phi_6_in1_valid, phi_6_in3_valid, phi_6_in2_valid}), .ready_in_bus({phi_6_in1_ready, phi_6_in3_ready, phi_6_in2_ready}), 
		.data_out_bus({phi_6_out1_data}), .valid_out_bus({phi_6_out1_valid}), .ready_out_bus({phi_6_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_7
		(.clk(phi_7_clk), .rst(phi_7_rst),
		.data_in_bus({{5'b0, phi_7_in1_data}, phi_7_in3_data, phi_7_in2_data}), .valid_in_bus({phi_7_in1_valid, phi_7_in3_valid, phi_7_in2_valid}), .ready_in_bus({phi_7_in1_ready, phi_7_in3_ready, phi_7_in2_ready}), 
		.data_out_bus({phi_7_out1_data}), .valid_out_bus({phi_7_out1_valid}), .ready_out_bus({phi_7_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_2
		(.clk(cst_2_clk), .rst(cst_2_rst),
		.data_in_bus({3'd5}), .valid_in_bus({cst_2_in1_valid}), .ready_in_bus({cst_2_in1_ready}), 
		.data_out_bus({cst_2_out1_data}), .valid_out_bus({cst_2_out1_valid}), .ready_out_bus({cst_2_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(11), .DATA_OUT_SIZE(11)) shl_op_shl_8
		(.clk(shl_8_clk), .rst(shl_8_rst),
		.data_in_bus({shl_8_in2_data, shl_8_in1_data}), .valid_in_bus({shl_8_in2_valid, shl_8_in1_valid}), .ready_in_bus({shl_8_in2_ready, shl_8_in1_ready}), 
		.data_out_bus({shl_8_out1_data}), .valid_out_bus({shl_8_out1_valid}), .ready_out_bus({shl_8_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(12), .DATA_OUT_SIZE(12)) add_op_add_9
		(.clk(add_9_clk), .rst(add_9_rst),
		.data_in_bus({add_9_in2_data, add_9_in1_data}), .valid_in_bus({add_9_in2_valid, add_9_in1_valid}), .ready_in_bus({add_9_in2_ready, add_9_in1_ready}), 
		.data_out_bus({add_9_out1_data}), .valid_out_bus({add_9_out1_valid}), .ready_out_bus({add_9_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(12), .DATA_SIZE(32)) mc_load_op_load_12
		(.clk(load_12_clk), .rst(load_12_rst),
		.data_in_bus({load_12_in1_data}), .address_in_bus({load_12_in2_data}), .valid_in_bus({load_12_in2_valid, load_12_in1_valid}), .ready_in_bus({load_12_in2_ready, load_12_in1_ready}), 
		.data_out_bus({load_12_out1_data}), .address_out_bus({load_12_out2_data}), .valid_out_bus({load_12_out2_valid, load_12_out1_valid}), .ready_out_bus({load_12_out2_ready, load_12_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_15
		(.clk(load_15_clk), .rst(load_15_rst),
		.data_in_bus({load_15_in1_data}), .address_in_bus({load_15_in2_data}), .valid_in_bus({load_15_in2_valid, load_15_in1_valid}), .ready_in_bus({load_15_in2_ready, load_15_in1_ready}), 
		.data_out_bus({load_15_out1_data}), .address_out_bus({load_15_out2_data}), .valid_out_bus({load_15_out2_valid, load_15_out1_valid}), .ready_out_bus({load_15_out2_ready, load_15_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_3
		(.clk(cst_3_clk), .rst(cst_3_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_3_in1_valid}), .ready_in_bus({cst_3_in1_ready}), 
		.data_out_bus({cst_3_out1_data}), .valid_out_bus({cst_3_out1_valid}), .ready_out_bus({cst_3_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_18
		(.clk(add_18_clk), .rst(add_18_rst),
		.data_in_bus({add_18_in2_data, add_18_in1_data}), .valid_in_bus({add_18_in2_valid, add_18_in1_valid}), .ready_in_bus({add_18_in2_ready, add_18_in1_ready}), 
		.data_out_bus({add_18_out1_data}), .valid_out_bus({add_18_out1_valid}), .ready_out_bus({add_18_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_4
		(.clk(cst_4_clk), .rst(cst_4_rst),
		.data_in_bus({6'd32}), .valid_in_bus({cst_4_in1_valid}), .ready_in_bus({cst_4_in1_ready}), 
		.data_out_bus({cst_4_out1_data}), .valid_out_bus({cst_4_out1_valid}), .ready_out_bus({cst_4_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_19
		(.clk(icmp_19_clk), .rst(icmp_19_rst),
		.data_in_bus({icmp_19_in2_data, icmp_19_in1_data}), .valid_in_bus({icmp_19_in2_valid, icmp_19_in1_valid}), .ready_in_bus({icmp_19_in2_ready, icmp_19_in1_ready}), 
		.data_out_bus({icmp_19_out1_data}), .valid_out_bus({icmp_19_out1_valid}), .ready_out_bus({icmp_19_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n2
		(.clk(phi_n2_clk), .rst(phi_n2_rst),
		.data_in_bus({phi_n2_in2_data, phi_n2_in1_data}), .valid_in_bus({phi_n2_in2_valid, phi_n2_in1_valid}), .ready_in_bus({phi_n2_in2_ready, phi_n2_in1_ready}), 
		.data_out_bus({phi_n2_out1_data}), .valid_out_bus({phi_n2_out1_valid}), .ready_out_bus({phi_n2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_1
		(.clk(fork_1_clk), .rst(fork_1_rst),
		.data_in_bus({fork_1_in1_data}), .valid_in_bus({fork_1_in1_valid}), .ready_in_bus({fork_1_in1_ready}), 
		.data_out_bus({fork_1_out3_data, fork_1_out2_data, fork_1_out1_data}), .valid_out_bus({fork_1_out3_valid, fork_1_out2_valid, fork_1_out1_valid}), .ready_out_bus({fork_1_out3_ready, fork_1_out2_ready, fork_1_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_3
		(.clk(fork_3_clk), .rst(fork_3_rst),
		.data_in_bus({fork_3_in1_data}), .valid_in_bus({fork_3_in1_valid}), .ready_in_bus({fork_3_in1_ready}), 
		.data_out_bus({fork_3_out2_data, fork_3_out1_data}), .valid_out_bus({fork_3_out2_valid, fork_3_out1_valid}), .ready_out_bus({fork_3_out2_ready, fork_3_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_11
		(.clk(fork_11_clk), .rst(fork_11_rst),
		.data_in_bus({fork_11_in1_data}), .valid_in_bus({fork_11_in1_valid}), .ready_in_bus({fork_11_in1_ready}), 
		.data_out_bus({fork_11_out2_data, fork_11_out1_data}), .valid_out_bus({fork_11_out2_valid, fork_11_out1_valid}), .ready_out_bus({fork_11_out2_ready, fork_11_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_4
		(.clk(branch_4_clk), .rst(branch_4_rst),
		.data_in_bus({{31'b0, branch_4_in2_data}, branch_4_in1_data}), .valid_in_bus({branch_4_in2_valid, branch_4_in1_valid}), .ready_in_bus({branch_4_in2_ready, branch_4_in1_ready}), 
		.data_out_bus({branch_4_out2_data, branch_4_out1_data}), .valid_out_bus({branch_4_out2_valid, branch_4_out1_valid}), .ready_out_bus({branch_4_out2_ready, branch_4_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_5
		(.clk(branch_5_clk), .rst(branch_5_rst),
		.data_in_bus({{5'b0, branch_5_in2_data}, branch_5_in1_data}), .valid_in_bus({branch_5_in2_valid, branch_5_in1_valid}), .ready_in_bus({branch_5_in2_ready, branch_5_in1_ready}), 
		.data_out_bus({branch_5_out2_data, branch_5_out1_data}), .valid_out_bus({branch_5_out2_valid, branch_5_out1_valid}), .ready_out_bus({branch_5_out2_ready, branch_5_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_6
		(.clk(branch_6_clk), .rst(branch_6_rst),
		.data_in_bus({{5'b0, branch_6_in2_data}, branch_6_in1_data}), .valid_in_bus({branch_6_in2_valid, branch_6_in1_valid}), .ready_in_bus({branch_6_in2_ready, branch_6_in1_ready}), 
		.data_out_bus({branch_6_out2_data, branch_6_out1_data}), .valid_out_bus({branch_6_out2_valid, branch_6_out1_valid}), .ready_out_bus({branch_6_out2_ready, branch_6_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_16
		(.clk(fork_16_clk), .rst(fork_16_rst),
		.data_in_bus({fork_16_in1_data}), .valid_in_bus({fork_16_in1_valid}), .ready_in_bus({fork_16_in1_ready}), 
		.data_out_bus({fork_16_out4_data, fork_16_out3_data, fork_16_out2_data, fork_16_out1_data}), .valid_out_bus({fork_16_out4_valid, fork_16_out3_valid, fork_16_out2_valid, fork_16_out1_valid}), .ready_out_bus({fork_16_out4_ready, fork_16_out3_ready, fork_16_out2_ready, fork_16_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_7
		(.clk(phiC_7_clk), .rst(phiC_7_rst),
		.data_in_bus({phiC_7_in2_data, phiC_7_in1_data}), .valid_in_bus({phiC_7_in2_valid, phiC_7_in1_valid}), .ready_in_bus({phiC_7_in2_ready, phiC_7_in1_ready}), 
		.data_out_bus({phiC_7_out2_data, phiC_7_out1_data}), .valid_out_bus({phiC_7_out2_valid, phiC_7_out1_valid}), .ready_out_bus({phiC_7_out2_ready, phiC_7_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_18
		(.clk(branchC_18_clk), .rst(branchC_18_rst),
		.data_in_bus({{branchC_18_in2_data}, branchC_18_in1_data}), .valid_in_bus({branchC_18_in2_valid, branchC_18_in1_valid}), .ready_in_bus({branchC_18_in2_ready, branchC_18_in1_ready}), 
		.data_out_bus({branchC_18_out2_data, branchC_18_out1_data}), .valid_out_bus({branchC_18_out2_valid, branchC_18_out1_valid}), .ready_out_bus({branchC_18_out2_ready, branchC_18_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_0
		(.clk(source_0_clk), .rst(source_0_rst),
		.data_out_bus({source_0_out1_data}), .valid_out_bus({source_0_out1_valid}), .ready_out_bus({source_0_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_1
		(.clk(source_1_clk), .rst(source_1_rst),
		.data_out_bus({source_1_out1_data}), .valid_out_bus({source_1_out1_valid}), .ready_out_bus({source_1_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_2
		(.clk(source_2_clk), .rst(source_2_rst),
		.data_out_bus({source_2_out1_data}), .valid_out_bus({source_2_out1_valid}), .ready_out_bus({source_2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_37
		(.clk(fork_37_clk), .rst(fork_37_rst),
		.data_in_bus({fork_37_in1_data}), .valid_in_bus({fork_37_in1_valid}), .ready_in_bus({fork_37_in1_ready}), 
		.data_out_bus({fork_37_out2_data, fork_37_out1_data}), .valid_out_bus({fork_37_out2_valid, fork_37_out1_valid}), .ready_out_bus({fork_37_out2_ready, fork_37_out1_ready}));

	mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_store_op_store_0
		(.clk(store_0_clk), .rst(store_0_rst),
		.data_in_bus({store_0_in1_data}), .address_in_bus({store_0_in2_data}), .valid_in_bus({store_0_in2_valid, store_0_in1_valid}), .ready_in_bus({store_0_in2_ready, store_0_in1_ready}), 
		.data_out_bus({store_0_out1_data}), .address_out_bus({store_0_out2_data}), .valid_out_bus({store_0_out2_valid, store_0_out1_valid}), .ready_out_bus({store_0_out2_ready, store_0_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_5
		(.clk(cst_5_clk), .rst(cst_5_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_5_in1_valid}), .ready_in_bus({cst_5_in1_ready}), 
		.data_out_bus({cst_5_out1_data}), .valid_out_bus({cst_5_out1_valid}), .ready_out_bus({cst_5_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_23
		(.clk(add_23_clk), .rst(add_23_rst),
		.data_in_bus({add_23_in2_data, add_23_in1_data}), .valid_in_bus({add_23_in2_valid, add_23_in1_valid}), .ready_in_bus({add_23_in2_ready, add_23_in1_ready}), 
		.data_out_bus({add_23_out1_data}), .valid_out_bus({add_23_out1_valid}), .ready_out_bus({add_23_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_6
		(.clk(cst_6_clk), .rst(cst_6_rst),
		.data_in_bus({6'd32}), .valid_in_bus({cst_6_in1_valid}), .ready_in_bus({cst_6_in1_ready}), 
		.data_out_bus({cst_6_out1_data}), .valid_out_bus({cst_6_out1_valid}), .ready_out_bus({cst_6_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_24
		(.clk(icmp_24_clk), .rst(icmp_24_rst),
		.data_in_bus({icmp_24_in2_data, icmp_24_in1_data}), .valid_in_bus({icmp_24_in2_valid, icmp_24_in1_valid}), .ready_in_bus({icmp_24_in2_ready, icmp_24_in1_ready}), 
		.data_out_bus({icmp_24_out1_data}), .valid_out_bus({icmp_24_out1_valid}), .ready_out_bus({icmp_24_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n0
		(.clk(phi_n0_clk), .rst(phi_n0_rst),
		.data_in_bus({phi_n0_in1_data}), .valid_in_bus({phi_n0_in1_valid}), .ready_in_bus({phi_n0_in1_ready}), 
		.data_out_bus({phi_n0_out1_data}), .valid_out_bus({phi_n0_out1_valid}), .ready_out_bus({phi_n0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n1
		(.clk(phi_n1_clk), .rst(phi_n1_rst),
		.data_in_bus({phi_n1_in1_data}), .valid_in_bus({phi_n1_in1_valid}), .ready_in_bus({phi_n1_in1_ready}), 
		.data_out_bus({phi_n1_out1_data}), .valid_out_bus({phi_n1_out1_valid}), .ready_out_bus({phi_n1_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_4
		(.clk(fork_4_clk), .rst(fork_4_rst),
		.data_in_bus({fork_4_in1_data}), .valid_in_bus({fork_4_in1_valid}), .ready_in_bus({fork_4_in1_ready}), 
		.data_out_bus({fork_4_out2_data, fork_4_out1_data}), .valid_out_bus({fork_4_out2_valid, fork_4_out1_valid}), .ready_out_bus({fork_4_out2_ready, fork_4_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_10
		(.clk(fork_10_clk), .rst(fork_10_rst),
		.data_in_bus({fork_10_in1_data}), .valid_in_bus({fork_10_in1_valid}), .ready_in_bus({fork_10_in1_ready}), 
		.data_out_bus({fork_10_out2_data, fork_10_out1_data}), .valid_out_bus({fork_10_out2_valid, fork_10_out1_valid}), .ready_out_bus({fork_10_out2_ready, fork_10_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_7
		(.clk(branch_7_clk), .rst(branch_7_rst),
		.data_in_bus({{5'b0, branch_7_in2_data}, branch_7_in1_data}), .valid_in_bus({branch_7_in2_valid, branch_7_in1_valid}), .ready_in_bus({branch_7_in2_ready, branch_7_in1_ready}), 
		.data_out_bus({branch_7_out2_data, branch_7_out1_data}), .valid_out_bus({branch_7_out2_valid, branch_7_out1_valid}), .ready_out_bus({branch_7_out2_ready, branch_7_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_14
		(.clk(cst_14_clk), .rst(cst_14_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_14_in1_valid}), .ready_in_bus({cst_14_in1_ready}), 
		.data_out_bus({cst_14_out1_data}), .valid_out_bus({cst_14_out1_valid}), .ready_out_bus({cst_14_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_8
		(.clk(phiC_8_clk), .rst(phiC_8_rst),
		.data_in_bus({phiC_8_in1_data}), .valid_in_bus({phiC_8_in1_valid}), .ready_in_bus({phiC_8_in1_ready}), 
		.data_out_bus({phiC_8_out1_data}), .valid_out_bus({phiC_8_out1_valid}), .ready_out_bus({phiC_8_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_27
		(.clk(forkC_27_clk), .rst(forkC_27_rst),
		.data_in_bus({forkC_27_in1_data}), .valid_in_bus({forkC_27_in1_valid}), .ready_in_bus({forkC_27_in1_ready}), 
		.data_out_bus({forkC_27_out2_data, forkC_27_out1_data}), .valid_out_bus({forkC_27_out2_valid, forkC_27_out1_valid}), .ready_out_bus({forkC_27_out2_ready, forkC_27_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_19
		(.clk(branchC_19_clk), .rst(branchC_19_rst),
		.data_in_bus({{branchC_19_in2_data}, branchC_19_in1_data}), .valid_in_bus({branchC_19_in2_valid, branchC_19_in1_valid}), .ready_in_bus({branchC_19_in2_ready, branchC_19_in1_ready}), 
		.data_out_bus({branchC_19_out2_data, branchC_19_out1_data}), .valid_out_bus({branchC_19_out2_valid, branchC_19_out1_valid}), .ready_out_bus({branchC_19_out2_ready, branchC_19_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_28
		(.clk(fork_28_clk), .rst(fork_28_rst),
		.data_in_bus({fork_28_in1_data}), .valid_in_bus({fork_28_in1_valid}), .ready_in_bus({fork_28_in1_ready}), 
		.data_out_bus({fork_28_out2_data, fork_28_out1_data}), .valid_out_bus({fork_28_out2_valid, fork_28_out1_valid}), .ready_out_bus({fork_28_out2_ready, fork_28_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_3
		(.clk(source_3_clk), .rst(source_3_rst),
		.data_out_bus({source_3_out1_data}), .valid_out_bus({source_3_out1_valid}), .ready_out_bus({source_3_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_4
		(.clk(source_4_clk), .rst(source_4_rst),
		.data_out_bus({source_4_out1_data}), .valid_out_bus({source_4_out1_valid}), .ready_out_bus({source_4_out1_ready}));

	ret_op #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) ret_op_ret_0
		(.clk(ret_0_clk), .rst(ret_0_rst),
		.data_in_bus({ret_0_in1_data}), .valid_in_bus({ret_0_in1_valid}), .ready_in_bus({ret_0_in1_ready}), 
		.data_out_bus({ret_0_out1_data}), .valid_out_bus({ret_0_out1_valid}), .ready_out_bus({ret_0_out1_ready}));

	end_node #(.INPUTS(1), .OUTPUTS(1), .MEMORY_INPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) end_node_end_0
		(.clk(end_0_clk), .rst(end_0_rst),
		.data_in_bus({end_0_in6_data}), .valid_in_bus({end_0_in6_valid}), .ready_in_bus({end_0_in6_ready}), .e_valid_bus({end_0_in5_valid, end_0_in4_valid, end_0_in3_valid, end_0_in2_valid, end_0_in1_valid}), .e_ready_bus({end_0_in5_ready, end_0_in4_ready, end_0_in3_ready, end_0_in2_ready, end_0_in1_ready}), 
		.data_out_bus({end_0_out1_data}), .valid_out_bus({end_0_out1_valid}), .ready_out_bus({end_0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_13
		(.clk(phiC_13_clk), .rst(phiC_13_rst),
		.data_in_bus({phiC_13_in1_data}), .valid_in_bus({phiC_13_in1_valid}), .ready_in_bus({phiC_13_in1_ready}), 
		.data_out_bus({phiC_13_out1_data}), .valid_out_bus({phiC_13_out1_valid}), .ready_out_bus({phiC_13_out1_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_x1
		(.clk(MC_x1_clk), .rst(MC_x1_rst),
		.io_storeDataOut(x1_dout0), .io_storeAddrOut(x1_address0), .io_storeEnable(x1_we0),
		.io_loadDataIn(x1_din1), .io_loadAddrOut(x1_address1), .io_loadEnable(x1_ce1),
		.io_bbpValids({MC_x1_in1_valid}), .io_bb_stCountArray({MC_x1_in1_data}), .io_bbReadyToPrevs({MC_x1_in1_ready}), .io_rdPortsPrev_ready({MC_x1_in2_ready}), .io_rdPortsPrev_valid({MC_x1_in2_valid}), .io_rdPortsPrev_bits({MC_x1_in2_data}), 	
	.io_wrAddrPorts_ready({MC_x1_in3_ready}), .io_wrAddrPorts_valid({MC_x1_in3_valid}), .io_wrAddrPorts_bits({MC_x1_in3_data}), 	
	.io_wrDataPorts_ready({MC_x1_in4_ready}), .io_wrDataPorts_valid({MC_x1_in4_valid}), .io_wrDataPorts_bits({MC_x1_in4_data}), 	
	.io_rdPortsNext_ready({MC_x1_out1_ready}), .io_rdPortsNext_valid({MC_x1_out1_valid}), .io_rdPortsNext_bits({MC_x1_out1_data}), 	
	.io_Empty_Valid({MC_x1_out2_valid}), .io_Empty_Ready({MC_x1_out2_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(12), .BB_COUNT(1), .LOAD_COUNT(2), .STORE_COUNT(1))MemCont_MC_A
		(.clk(MC_A_clk), .rst(MC_A_rst),
		.io_storeDataOut(A_dout0), .io_storeAddrOut(A_address0), .io_storeEnable(A_we0),
		.io_loadDataIn(A_din1), .io_loadAddrOut(A_address1), .io_loadEnable(A_ce1),
		.io_bbpValids({MC_A_in3_valid}), .io_bb_stCountArray({MC_A_in3_data}), .io_bbReadyToPrevs({MC_A_in3_ready}), .io_rdPortsPrev_ready({MC_A_in2_ready, MC_A_in1_ready}), .io_rdPortsPrev_valid({MC_A_in2_valid, MC_A_in1_valid}), .io_rdPortsPrev_bits({MC_A_in2_data, MC_A_in1_data}), 	
	.io_wrAddrPorts_ready({MC_A_in4_ready}), .io_wrAddrPorts_valid({MC_A_in4_valid}), .io_wrAddrPorts_bits({MC_A_in4_data}), 	
	.io_wrDataPorts_ready({MC_A_in5_ready}), .io_wrDataPorts_valid({MC_A_in5_valid}), .io_wrDataPorts_bits({MC_A_in5_data}), 	
	.io_rdPortsNext_ready({MC_A_out2_ready, MC_A_out1_ready}), .io_rdPortsNext_valid({MC_A_out2_valid, MC_A_out1_valid}), .io_rdPortsNext_bits({MC_A_out2_data, MC_A_out1_data}), 	
	.io_Empty_Valid({MC_A_out3_valid}), .io_Empty_Ready({MC_A_out3_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_y1
		(.clk(MC_y1_clk), .rst(MC_y1_rst),
		.io_storeDataOut(y1_dout0), .io_storeAddrOut(y1_address0), .io_storeEnable(y1_we0),
		.io_loadDataIn(y1_din1), .io_loadAddrOut(y1_address1), .io_loadEnable(y1_ce1),
		.io_bbpValids({MC_y1_in2_valid}), .io_bb_stCountArray({MC_y1_in2_data}), .io_bbReadyToPrevs({MC_y1_in2_ready}), .io_rdPortsPrev_ready({MC_y1_in1_ready}), .io_rdPortsPrev_valid({MC_y1_in1_valid}), .io_rdPortsPrev_bits({MC_y1_in1_data}), 	
	.io_wrAddrPorts_ready({MC_y1_in3_ready}), .io_wrAddrPorts_valid({MC_y1_in3_valid}), .io_wrAddrPorts_bits({MC_y1_in3_data}), 	
	.io_wrDataPorts_ready({MC_y1_in4_ready}), .io_wrDataPorts_valid({MC_y1_in4_valid}), .io_wrDataPorts_bits({MC_y1_in4_data}), 	
	.io_rdPortsNext_ready({MC_y1_out1_ready}), .io_rdPortsNext_valid({MC_y1_out1_valid}), .io_rdPortsNext_bits({MC_y1_out1_data}), 	
	.io_Empty_Valid({MC_y1_out2_valid}), .io_Empty_Ready({MC_y1_out2_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_x2
		(.clk(MC_x2_clk), .rst(MC_x2_rst),
		.io_storeDataOut(x2_dout0), .io_storeAddrOut(x2_address0), .io_storeEnable(x2_we0),
		.io_loadDataIn(x2_din1), .io_loadAddrOut(x2_address1), .io_loadEnable(x2_ce1),
		.io_bbpValids({MC_x2_in1_valid}), .io_bb_stCountArray({MC_x2_in1_data}), .io_bbReadyToPrevs({MC_x2_in1_ready}), .io_rdPortsPrev_ready({MC_x2_in2_ready}), .io_rdPortsPrev_valid({MC_x2_in2_valid}), .io_rdPortsPrev_bits({MC_x2_in2_data}), 	
	.io_wrAddrPorts_ready({MC_x2_in3_ready}), .io_wrAddrPorts_valid({MC_x2_in3_valid}), .io_wrAddrPorts_bits({MC_x2_in3_data}), 	
	.io_wrDataPorts_ready({MC_x2_in4_ready}), .io_wrDataPorts_valid({MC_x2_in4_valid}), .io_wrDataPorts_bits({MC_x2_in4_data}), 	
	.io_rdPortsNext_ready({MC_x2_out1_ready}), .io_rdPortsNext_valid({MC_x2_out1_valid}), .io_rdPortsNext_bits({MC_x2_out1_data}), 	
	.io_Empty_Valid({MC_x2_out2_valid}), .io_Empty_Ready({MC_x2_out2_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_y2
		(.clk(MC_y2_clk), .rst(MC_y2_rst),
		.io_storeDataOut(y2_dout0), .io_storeAddrOut(y2_address0), .io_storeEnable(y2_we0),
		.io_loadDataIn(y2_din1), .io_loadAddrOut(y2_address1), .io_loadEnable(y2_ce1),
		.io_bbpValids({MC_y2_in2_valid}), .io_bb_stCountArray({MC_y2_in2_data}), .io_bbReadyToPrevs({MC_y2_in2_ready}), .io_rdPortsPrev_ready({MC_y2_in1_ready}), .io_rdPortsPrev_valid({MC_y2_in1_valid}), .io_rdPortsPrev_bits({MC_y2_in1_data}), 	
	.io_wrAddrPorts_ready({MC_y2_in3_ready}), .io_wrAddrPorts_valid({MC_y2_in3_valid}), .io_wrAddrPorts_bits({MC_y2_in3_data}), 	
	.io_wrDataPorts_ready({MC_y2_in4_ready}), .io_wrDataPorts_valid({MC_y2_in4_valid}), .io_wrDataPorts_bits({MC_y2_in4_data}), 	
	.io_rdPortsNext_ready({MC_y2_out1_ready}), .io_rdPortsNext_valid({MC_y2_out1_valid}), .io_rdPortsNext_bits({MC_y2_out1_data}), 	
	.io_Empty_Valid({MC_y2_out2_valid}), .io_Empty_Ready({MC_y2_out2_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_0
		(.clk(sink_0_clk), .rst(sink_0_rst),
		.data_in_bus({sink_0_in1_data}), .valid_in_bus({sink_0_in1_valid}), .ready_in_bus({sink_0_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_1
		(.clk(sink_1_clk), .rst(sink_1_rst),
		.data_in_bus({sink_1_in1_data}), .valid_in_bus({sink_1_in1_valid}), .ready_in_bus({sink_1_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_2
		(.clk(sink_2_clk), .rst(sink_2_rst),
		.data_in_bus({sink_2_in1_data}), .valid_in_bus({sink_2_in1_valid}), .ready_in_bus({sink_2_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_3
		(.clk(sink_3_clk), .rst(sink_3_rst),
		.data_in_bus({sink_3_in1_data}), .valid_in_bus({sink_3_in1_valid}), .ready_in_bus({sink_3_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_4
		(.clk(sink_4_clk), .rst(sink_4_rst),
		.data_in_bus({sink_4_in1_data}), .valid_in_bus({sink_4_in1_valid}), .ready_in_bus({sink_4_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_5
		(.clk(sink_5_clk), .rst(sink_5_rst),
		.data_in_bus({sink_5_in1_data}), .valid_in_bus({sink_5_in1_valid}), .ready_in_bus({sink_5_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_6
		(.clk(sink_6_clk), .rst(sink_6_rst),
		.data_in_bus({sink_6_in1_data}), .valid_in_bus({sink_6_in1_valid}), .ready_in_bus({sink_6_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_7
		(.clk(sink_7_clk), .rst(sink_7_rst),
		.data_in_bus({sink_7_in1_data}), .valid_in_bus({sink_7_in1_valid}), .ready_in_bus({sink_7_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_8
		(.clk(sink_8_clk), .rst(sink_8_rst),
		.data_in_bus({sink_8_in1_data}), .valid_in_bus({sink_8_in1_valid}), .ready_in_bus({sink_8_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_9
		(.clk(sink_9_clk), .rst(sink_9_rst),
		.data_in_bus({sink_9_in1_data}), .valid_in_bus({sink_9_in1_valid}), .ready_in_bus({sink_9_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_10
		(.clk(sink_10_clk), .rst(sink_10_rst),
		.data_in_bus({sink_10_in1_data}), .valid_in_bus({sink_10_in1_valid}), .ready_in_bus({sink_10_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_11
		(.clk(sink_11_clk), .rst(sink_11_rst),
		.data_in_bus({sink_11_in1_data}), .valid_in_bus({sink_11_in1_valid}), .ready_in_bus({sink_11_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_12
		(.clk(sink_12_clk), .rst(sink_12_rst),
		.data_in_bus({sink_12_in1_data}), .valid_in_bus({sink_12_in1_valid}), .ready_in_bus({sink_12_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_13
		(.clk(sink_13_clk), .rst(sink_13_rst),
		.data_in_bus({sink_13_in1_data}), .valid_in_bus({sink_13_in1_valid}), .ready_in_bus({sink_13_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_14
		(.clk(sink_14_clk), .rst(sink_14_rst),
		.data_in_bus({sink_14_in1_data}), .valid_in_bus({sink_14_in1_valid}), .ready_in_bus({sink_14_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_15
		(.clk(sink_15_clk), .rst(sink_15_rst),
		.data_in_bus({sink_15_in1_data}), .valid_in_bus({sink_15_in1_valid}), .ready_in_bus({sink_15_in1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_100
		(.clk(Buffer_100_clk), .rst(Buffer_100_rst),
		.data_in_bus({Buffer_100_in1_data}), .valid_in_bus({Buffer_100_in1_valid}), .ready_in_bus({Buffer_100_in1_ready}), 
		.data_out_bus({Buffer_100_out1_data}), .valid_out_bus({Buffer_100_out1_valid}), .ready_out_bus({Buffer_100_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_101
		(.clk(Buffer_101_clk), .rst(Buffer_101_rst),
		.data_in_bus({Buffer_101_in1_data}), .valid_in_bus({Buffer_101_in1_valid}), .ready_in_bus({Buffer_101_in1_ready}), 
		.data_out_bus({Buffer_101_out1_data}), .valid_out_bus({Buffer_101_out1_valid}), .ready_out_bus({Buffer_101_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_102
		(.clk(Buffer_102_clk), .rst(Buffer_102_rst),
		.data_in_bus({Buffer_102_in1_data}), .valid_in_bus({Buffer_102_in1_valid}), .ready_in_bus({Buffer_102_in1_ready}), 
		.data_out_bus({Buffer_102_out1_data}), .valid_out_bus({Buffer_102_out1_valid}), .ready_out_bus({Buffer_102_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_103
		(.clk(Buffer_103_clk), .rst(Buffer_103_rst),
		.data_in_bus({Buffer_103_in1_data}), .valid_in_bus({Buffer_103_in1_valid}), .ready_in_bus({Buffer_103_in1_ready}), 
		.data_out_bus({Buffer_103_out1_data}), .valid_out_bus({Buffer_103_out1_valid}), .ready_out_bus({Buffer_103_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_104
		(.clk(Buffer_104_clk), .rst(Buffer_104_rst),
		.data_in_bus({Buffer_104_in1_data}), .valid_in_bus({Buffer_104_in1_valid}), .ready_in_bus({Buffer_104_in1_ready}), 
		.data_out_bus({Buffer_104_out1_data}), .valid_out_bus({Buffer_104_out1_valid}), .ready_out_bus({Buffer_104_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_105
		(.clk(Buffer_105_clk), .rst(Buffer_105_rst),
		.data_in_bus({Buffer_105_in1_data}), .valid_in_bus({Buffer_105_in1_valid}), .ready_in_bus({Buffer_105_in1_ready}), 
		.data_out_bus({Buffer_105_out1_data}), .valid_out_bus({Buffer_105_out1_valid}), .ready_out_bus({Buffer_105_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_106
		(.clk(Buffer_106_clk), .rst(Buffer_106_rst),
		.data_in_bus({Buffer_106_in1_data}), .valid_in_bus({Buffer_106_in1_valid}), .ready_in_bus({Buffer_106_in1_ready}), 
		.data_out_bus({Buffer_106_out1_data}), .valid_out_bus({Buffer_106_out1_valid}), .ready_out_bus({Buffer_106_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_107
		(.clk(Buffer_107_clk), .rst(Buffer_107_rst),
		.data_in_bus({Buffer_107_in1_data}), .valid_in_bus({Buffer_107_in1_valid}), .ready_in_bus({Buffer_107_in1_ready}), 
		.data_out_bus({Buffer_107_out1_data}), .valid_out_bus({Buffer_107_out1_valid}), .ready_out_bus({Buffer_107_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_108
		(.clk(Buffer_108_clk), .rst(Buffer_108_rst),
		.data_in_bus({Buffer_108_in1_data}), .valid_in_bus({Buffer_108_in1_valid}), .ready_in_bus({Buffer_108_in1_ready}), 
		.data_out_bus({Buffer_108_out1_data}), .valid_out_bus({Buffer_108_out1_valid}), .ready_out_bus({Buffer_108_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_109
		(.clk(Buffer_109_clk), .rst(Buffer_109_rst),
		.data_in_bus({Buffer_109_in1_data}), .valid_in_bus({Buffer_109_in1_valid}), .ready_in_bus({Buffer_109_in1_ready}), 
		.data_out_bus({Buffer_109_out1_data}), .valid_out_bus({Buffer_109_out1_valid}), .ready_out_bus({Buffer_109_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_110
		(.clk(Buffer_110_clk), .rst(Buffer_110_rst),
		.data_in_bus({Buffer_110_in1_data}), .valid_in_bus({Buffer_110_in1_valid}), .ready_in_bus({Buffer_110_in1_ready}), 
		.data_out_bus({Buffer_110_out1_data}), .valid_out_bus({Buffer_110_out1_valid}), .ready_out_bus({Buffer_110_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_111
		(.clk(Buffer_111_clk), .rst(Buffer_111_rst),
		.data_in_bus({Buffer_111_in1_data}), .valid_in_bus({Buffer_111_in1_valid}), .ready_in_bus({Buffer_111_in1_ready}), 
		.data_out_bus({Buffer_111_out1_data}), .valid_out_bus({Buffer_111_out1_valid}), .ready_out_bus({Buffer_111_out1_ready}));

	and_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) and_op_and_300
		(.clk(and_300_clk), .rst(and_300_rst),
		.data_in_bus({and_300_in2_data, and_300_in1_data}), .valid_in_bus({and_300_in2_valid, and_300_in1_valid}), .ready_in_bus({and_300_in2_ready, and_300_in1_ready}), 
		.data_out_bus({and_300_out1_data}), .valid_out_bus({and_300_out1_valid}), .ready_out_bus({and_300_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_300
		(.clk(Buffer_300_clk), .rst(Buffer_300_rst),
		.data_in_bus({Buffer_300_in1_data}), .valid_in_bus({Buffer_300_in1_valid}), .ready_in_bus({Buffer_300_in1_ready}), 
		.data_out_bus({Buffer_300_out1_data}), .valid_out_bus({Buffer_300_out1_valid}), .ready_out_bus({Buffer_300_out1_ready}));

	and_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) and_op_and_301
		(.clk(and_301_clk), .rst(and_301_rst),
		.data_in_bus({and_301_in2_data, and_301_in1_data}), .valid_in_bus({and_301_in2_valid, and_301_in1_valid}), .ready_in_bus({and_301_in2_ready, and_301_in1_ready}), 
		.data_out_bus({and_301_out1_data}), .valid_out_bus({and_301_out1_valid}), .ready_out_bus({and_301_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_301
		(.clk(Buffer_301_clk), .rst(Buffer_301_rst),
		.data_in_bus({Buffer_301_in1_data}), .valid_in_bus({Buffer_301_in1_valid}), .ready_in_bus({Buffer_301_in1_ready}), 
		.data_out_bus({Buffer_301_out1_data}), .valid_out_bus({Buffer_301_out1_valid}), .ready_out_bus({Buffer_301_out1_ready}));

	and_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) and_op_and_302
		(.clk(and_302_clk), .rst(and_302_rst),
		.data_in_bus({and_302_in2_data, and_302_in1_data}), .valid_in_bus({and_302_in2_valid, and_302_in1_valid}), .ready_in_bus({and_302_in2_ready, and_302_in1_ready}), 
		.data_out_bus({and_302_out1_data}), .valid_out_bus({and_302_out1_valid}), .ready_out_bus({and_302_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_302
		(.clk(Buffer_302_clk), .rst(Buffer_302_rst),
		.data_in_bus({Buffer_302_in1_data}), .valid_in_bus({Buffer_302_in1_valid}), .ready_in_bus({Buffer_302_in1_ready}), 
		.data_out_bus({Buffer_302_out1_data}), .valid_out_bus({Buffer_302_out1_valid}), .ready_out_bus({Buffer_302_out1_ready}));

	and_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) and_op_and_303
		(.clk(and_303_clk), .rst(and_303_rst),
		.data_in_bus({and_303_in2_data, and_303_in1_data}), .valid_in_bus({and_303_in2_valid, and_303_in1_valid}), .ready_in_bus({and_303_in2_ready, and_303_in1_ready}), 
		.data_out_bus({and_303_out1_data}), .valid_out_bus({and_303_out1_valid}), .ready_out_bus({and_303_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_303
		(.clk(Buffer_303_clk), .rst(Buffer_303_rst),
		.data_in_bus({Buffer_303_in1_data}), .valid_in_bus({Buffer_303_in1_valid}), .ready_in_bus({Buffer_303_in1_ready}), 
		.data_out_bus({Buffer_303_out1_data}), .valid_out_bus({Buffer_303_out1_valid}), .ready_out_bus({Buffer_303_out1_ready}));

endmodule

