module gaussian(
	input clk,
	input rst,

	input [0 : 0]start_in,
	input start_valid,
	output start_ready,

	output [0 : 0]end_out,
	output end_valid,
	input end_ready,

	output [9 : 0]A_address0,
	output A_ce0,
	output A_we0,
	output [31 : 0]A_dout0,
	input [31 : 0]A_din0,
	output [9 : 0]A_address1,
	output A_ce1,
	output A_we1,
	output [31 : 0]A_dout1,
	input [31 : 0]A_din1,

	output [4 : 0]c_address0,
	output c_ce0,
	output c_we0,
	output [31 : 0]c_dout0,
	input [31 : 0]c_din0,
	output [4 : 0]c_address1,
	output c_ce1,
	output c_we1,
	output [31 : 0]c_dout1,
	input [31 : 0]c_din1

);

	wire brCst_block1_clk;
	wire brCst_block1_rst;
	wire [0 : 0]brCst_block1_in1_data;
	wire brCst_block1_in1_ready;
	wire brCst_block1_in1_valid;
	wire [0 : 0]brCst_block1_out1_data;
	wire brCst_block1_out1_ready;
	wire brCst_block1_out1_valid;

	wire cst_0_clk;
	wire cst_0_rst;
	wire [0 : 0]cst_0_in1_data;
	wire cst_0_in1_ready;
	wire cst_0_in1_valid;
	wire [0 : 0]cst_0_out1_data;
	wire cst_0_out1_ready;
	wire cst_0_out1_valid;

	wire branch_0_clk;
	wire branch_0_rst;
	wire [0 : 0]branch_0_in1_data;
	wire branch_0_in1_ready;
	wire branch_0_in1_valid;
	wire [0 : 0]branch_0_in2_data;
	wire branch_0_in2_ready;
	wire branch_0_in2_valid;
	wire [0 : 0]branch_0_out1_data;
	wire branch_0_out1_ready;
	wire branch_0_out1_valid;
	wire [0 : 0]branch_0_out2_data;
	wire branch_0_out2_ready;
	wire branch_0_out2_valid;

	wire start_0_clk;
	wire start_0_rst;
	wire [0 : 0]start_0_in1_data;
	wire start_0_in1_ready;
	wire start_0_in1_valid;
	wire [0 : 0]start_0_out1_data;
	wire start_0_out1_ready;
	wire start_0_out1_valid;

	wire forkC_17_clk;
	wire forkC_17_rst;
	wire [0 : 0]forkC_17_in1_data;
	wire forkC_17_in1_ready;
	wire forkC_17_in1_valid;
	wire [0 : 0]forkC_17_out1_data;
	wire forkC_17_out1_ready;
	wire forkC_17_out1_valid;
	wire [0 : 0]forkC_17_out2_data;
	wire forkC_17_out2_ready;
	wire forkC_17_out2_valid;
	wire [0 : 0]forkC_17_out3_data;
	wire forkC_17_out3_ready;
	wire forkC_17_out3_valid;

	wire branchC_14_clk;
	wire branchC_14_rst;
	wire [0 : 0]branchC_14_in1_data;
	wire branchC_14_in1_ready;
	wire branchC_14_in1_valid;
	wire [0 : 0]branchC_14_in2_data;
	wire branchC_14_in2_ready;
	wire branchC_14_in2_valid;
	wire [0 : 0]branchC_14_out1_data;
	wire branchC_14_out1_ready;
	wire branchC_14_out1_valid;
	wire [0 : 0]branchC_14_out2_data;
	wire branchC_14_out2_ready;
	wire branchC_14_out2_valid;

	wire fork_18_clk;
	wire fork_18_rst;
	wire [0 : 0]fork_18_in1_data;
	wire fork_18_in1_ready;
	wire fork_18_in1_valid;
	wire [0 : 0]fork_18_out1_data;
	wire fork_18_out1_ready;
	wire fork_18_out1_valid;
	wire [0 : 0]fork_18_out2_data;
	wire fork_18_out2_ready;
	wire fork_18_out2_valid;

	wire brCst_block3_clk;
	wire brCst_block3_rst;
	wire [0 : 0]brCst_block3_in1_data;
	wire brCst_block3_in1_ready;
	wire brCst_block3_in1_valid;
	wire [0 : 0]brCst_block3_out1_data;
	wire brCst_block3_out1_ready;
	wire brCst_block3_out1_valid;

	wire phi_n1_clk;
	wire phi_n1_rst;
	wire [5 : 0]phi_n1_in1_data;
	wire phi_n1_in1_ready;
	wire phi_n1_in1_valid;
	wire [5 : 0]phi_n1_out1_data;
	wire phi_n1_out1_ready;
	wire phi_n1_out1_valid;

	wire phi_n2_clk;
	wire phi_n2_rst;
	wire [4 : 0]phi_n2_in1_data;
	wire phi_n2_in1_ready;
	wire phi_n2_in1_valid;
	wire [4 : 0]phi_n2_out1_data;
	wire phi_n2_out1_ready;
	wire phi_n2_out1_valid;

	wire branch_3_clk;
	wire branch_3_rst;
	wire [5 : 0]branch_3_in1_data;
	wire branch_3_in1_ready;
	wire branch_3_in1_valid;
	wire [0 : 0]branch_3_in2_data;
	wire branch_3_in2_ready;
	wire branch_3_in2_valid;
	wire [5 : 0]branch_3_out1_data;
	wire branch_3_out1_ready;
	wire branch_3_out1_valid;
	wire [5 : 0]branch_3_out2_data;
	wire branch_3_out2_ready;
	wire branch_3_out2_valid;

	wire branch_4_clk;
	wire branch_4_rst;
	wire [4 : 0]branch_4_in1_data;
	wire branch_4_in1_ready;
	wire branch_4_in1_valid;
	wire [0 : 0]branch_4_in2_data;
	wire branch_4_in2_ready;
	wire branch_4_in2_valid;
	wire [4 : 0]branch_4_out1_data;
	wire branch_4_out1_ready;
	wire branch_4_out1_valid;
	wire [4 : 0]branch_4_out2_data;
	wire branch_4_out2_ready;
	wire branch_4_out2_valid;

	wire fork_11_clk;
	wire fork_11_rst;
	wire [0 : 0]fork_11_in1_data;
	wire fork_11_in1_ready;
	wire fork_11_in1_valid;
	wire [0 : 0]fork_11_out1_data;
	wire fork_11_out1_ready;
	wire fork_11_out1_valid;
	wire [0 : 0]fork_11_out2_data;
	wire fork_11_out2_ready;
	wire fork_11_out2_valid;
	wire [0 : 0]fork_11_out3_data;
	wire fork_11_out3_ready;
	wire fork_11_out3_valid;

	wire phiC_9_clk;
	wire phiC_9_rst;
	wire [0 : 0]phiC_9_in1_data;
	wire phiC_9_in1_ready;
	wire phiC_9_in1_valid;
	wire [0 : 0]phiC_9_out1_data;
	wire phiC_9_out1_ready;
	wire phiC_9_out1_valid;

	wire forkC_20_clk;
	wire forkC_20_rst;
	wire [0 : 0]forkC_20_in1_data;
	wire forkC_20_in1_ready;
	wire forkC_20_in1_valid;
	wire [0 : 0]forkC_20_out1_data;
	wire forkC_20_out1_ready;
	wire forkC_20_out1_valid;
	wire [0 : 0]forkC_20_out2_data;
	wire forkC_20_out2_ready;
	wire forkC_20_out2_valid;

	wire branchC_16_clk;
	wire branchC_16_rst;
	wire [0 : 0]branchC_16_in1_data;
	wire branchC_16_in1_ready;
	wire branchC_16_in1_valid;
	wire [0 : 0]branchC_16_in2_data;
	wire branchC_16_in2_ready;
	wire branchC_16_in2_valid;
	wire [0 : 0]branchC_16_out1_data;
	wire branchC_16_out1_ready;
	wire branchC_16_out1_valid;
	wire [0 : 0]branchC_16_out2_data;
	wire branchC_16_out2_ready;
	wire branchC_16_out2_valid;

	wire cst_9_clk;
	wire cst_9_rst;
	wire [0 : 0]cst_9_in1_data;
	wire cst_9_in1_ready;
	wire cst_9_in1_valid;
	wire [0 : 0]cst_9_out1_data;
	wire cst_9_out1_ready;
	wire cst_9_out1_valid;

	wire add_31_clk;
	wire add_31_rst;
	wire [4 : 0]add_31_in1_data;
	wire add_31_in1_ready;
	wire add_31_in1_valid;
	wire [4 : 0]add_31_in2_data;
	wire add_31_in2_ready;
	wire add_31_in2_valid;
	wire [4 : 0]add_31_out1_data;
	wire add_31_out1_ready;
	wire add_31_out1_valid;

	wire cst_10_clk;
	wire cst_10_rst;
	wire [3 : 0]cst_10_in1_data;
	wire cst_10_in1_ready;
	wire cst_10_in1_valid;
	wire [3 : 0]cst_10_out1_data;
	wire cst_10_out1_ready;
	wire cst_10_out1_valid;

	wire icmp_32_clk;
	wire icmp_32_rst;
	wire [5 : 0]icmp_32_in1_data;
	wire icmp_32_in1_ready;
	wire icmp_32_in1_valid;
	wire [5 : 0]icmp_32_in2_data;
	wire icmp_32_in2_ready;
	wire icmp_32_in2_valid;
	wire [0 : 0]icmp_32_out1_data;
	wire icmp_32_out1_ready;
	wire icmp_32_out1_valid;

	wire phi_n4_clk;
	wire phi_n4_rst;
	wire [4 : 0]phi_n4_in1_data;
	wire phi_n4_in1_ready;
	wire phi_n4_in1_valid;
	wire [4 : 0]phi_n4_out1_data;
	wire phi_n4_out1_ready;
	wire phi_n4_out1_valid;

	wire phi_n5_clk;
	wire phi_n5_rst;
	wire [4 : 0]phi_n5_in1_data;
	wire phi_n5_in1_ready;
	wire phi_n5_in1_valid;
	wire [4 : 0]phi_n5_out1_data;
	wire phi_n5_out1_ready;
	wire phi_n5_out1_valid;

	wire fork_5_clk;
	wire fork_5_rst;
	wire [4 : 0]fork_5_in1_data;
	wire fork_5_in1_ready;
	wire fork_5_in1_valid;
	wire [4 : 0]fork_5_out1_data;
	wire fork_5_out1_ready;
	wire fork_5_out1_valid;
	wire [4 : 0]fork_5_out2_data;
	wire fork_5_out2_ready;
	wire fork_5_out2_valid;

	wire branch_11_clk;
	wire branch_11_rst;
	wire [4 : 0]branch_11_in1_data;
	wire branch_11_in1_ready;
	wire branch_11_in1_valid;
	wire [0 : 0]branch_11_in2_data;
	wire branch_11_in2_ready;
	wire branch_11_in2_valid;
	wire [4 : 0]branch_11_out1_data;
	wire branch_11_out1_ready;
	wire branch_11_out1_valid;
	wire [4 : 0]branch_11_out2_data;
	wire branch_11_out2_ready;
	wire branch_11_out2_valid;

	wire branch_12_clk;
	wire branch_12_rst;
	wire [4 : 0]branch_12_in1_data;
	wire branch_12_in1_ready;
	wire branch_12_in1_valid;
	wire [0 : 0]branch_12_in2_data;
	wire branch_12_in2_ready;
	wire branch_12_in2_valid;
	wire [4 : 0]branch_12_out1_data;
	wire branch_12_out1_ready;
	wire branch_12_out1_valid;
	wire [4 : 0]branch_12_out2_data;
	wire branch_12_out2_ready;
	wire branch_12_out2_valid;

	wire fork_14_clk;
	wire fork_14_rst;
	wire [0 : 0]fork_14_in1_data;
	wire fork_14_in1_ready;
	wire fork_14_in1_valid;
	wire [0 : 0]fork_14_out1_data;
	wire fork_14_out1_ready;
	wire fork_14_out1_valid;
	wire [0 : 0]fork_14_out2_data;
	wire fork_14_out2_ready;
	wire fork_14_out2_valid;
	wire [0 : 0]fork_14_out3_data;
	wire fork_14_out3_ready;
	wire fork_14_out3_valid;

	wire phiC_12_clk;
	wire phiC_12_rst;
	wire [0 : 0]phiC_12_in1_data;
	wire phiC_12_in1_ready;
	wire phiC_12_in1_valid;
	wire [0 : 0]phiC_12_out1_data;
	wire phiC_12_out1_ready;
	wire phiC_12_out1_valid;

	wire branchC_19_clk;
	wire branchC_19_rst;
	wire [0 : 0]branchC_19_in1_data;
	wire branchC_19_in1_ready;
	wire branchC_19_in1_valid;
	wire [0 : 0]branchC_19_in2_data;
	wire branchC_19_in2_ready;
	wire branchC_19_in2_valid;
	wire [0 : 0]branchC_19_out1_data;
	wire branchC_19_out1_ready;
	wire branchC_19_out1_valid;
	wire [0 : 0]branchC_19_out2_data;
	wire branchC_19_out2_ready;
	wire branchC_19_out2_valid;

	wire source_7_clk;
	wire source_7_rst;
	wire [0 : 0]source_7_out1_data;
	wire source_7_out1_ready;
	wire source_7_out1_valid;

	wire source_8_clk;
	wire source_8_rst;
	wire [3 : 0]source_8_out1_data;
	wire source_8_out1_ready;
	wire source_8_out1_valid;

	wire cst_11_clk;
	wire cst_11_rst;
	wire [0 : 0]cst_11_in1_data;
	wire cst_11_in1_ready;
	wire cst_11_in1_valid;
	wire [0 : 0]cst_11_out1_data;
	wire cst_11_out1_ready;
	wire cst_11_out1_valid;

	wire add_34_clk;
	wire add_34_rst;
	wire [4 : 0]add_34_in1_data;
	wire add_34_in1_ready;
	wire add_34_in1_valid;
	wire [4 : 0]add_34_in2_data;
	wire add_34_in2_ready;
	wire add_34_in2_valid;
	wire [4 : 0]add_34_out1_data;
	wire add_34_out1_ready;
	wire add_34_out1_valid;

	wire cst_12_clk;
	wire cst_12_rst;
	wire [4 : 0]cst_12_in1_data;
	wire cst_12_in1_ready;
	wire cst_12_in1_valid;
	wire [4 : 0]cst_12_out1_data;
	wire cst_12_out1_ready;
	wire cst_12_out1_valid;

	wire icmp_35_clk;
	wire icmp_35_rst;
	wire [4 : 0]icmp_35_in1_data;
	wire icmp_35_in1_ready;
	wire icmp_35_in1_valid;
	wire [4 : 0]icmp_35_in2_data;
	wire icmp_35_in2_ready;
	wire icmp_35_in2_valid;
	wire [0 : 0]icmp_35_out1_data;
	wire icmp_35_out1_ready;
	wire icmp_35_out1_valid;

	wire phi_n0_clk;
	wire phi_n0_rst;
	wire [4 : 0]phi_n0_in1_data;
	wire phi_n0_in1_ready;
	wire phi_n0_in1_valid;
	wire [4 : 0]phi_n0_in2_data;
	wire phi_n0_in2_ready;
	wire phi_n0_in2_valid;
	wire [4 : 0]phi_n0_out1_data;
	wire phi_n0_out1_ready;
	wire phi_n0_out1_valid;

	wire fork_4_clk;
	wire fork_4_rst;
	wire [4 : 0]fork_4_in1_data;
	wire fork_4_in1_ready;
	wire fork_4_in1_valid;
	wire [4 : 0]fork_4_out1_data;
	wire fork_4_out1_ready;
	wire fork_4_out1_valid;
	wire [4 : 0]fork_4_out2_data;
	wire fork_4_out2_ready;
	wire fork_4_out2_valid;

	wire branch_13_clk;
	wire branch_13_rst;
	wire [4 : 0]branch_13_in1_data;
	wire branch_13_in1_ready;
	wire branch_13_in1_valid;
	wire [0 : 0]branch_13_in2_data;
	wire branch_13_in2_ready;
	wire branch_13_in2_valid;
	wire [4 : 0]branch_13_out1_data;
	wire branch_13_out1_ready;
	wire branch_13_out1_valid;
	wire [4 : 0]branch_13_out2_data;
	wire branch_13_out2_ready;
	wire branch_13_out2_valid;

	wire phiC_13_clk;
	wire phiC_13_rst;
	wire [0 : 0]phiC_13_in1_data;
	wire phiC_13_in1_ready;
	wire phiC_13_in1_valid;
	wire [0 : 0]phiC_13_in2_data;
	wire phiC_13_in2_ready;
	wire phiC_13_in2_valid;
	wire [0 : 0]phiC_13_out1_data;
	wire phiC_13_out1_ready;
	wire phiC_13_out1_valid;

	wire branchC_20_clk;
	wire branchC_20_rst;
	wire [0 : 0]branchC_20_in1_data;
	wire branchC_20_in1_ready;
	wire branchC_20_in1_valid;
	wire [0 : 0]branchC_20_in2_data;
	wire branchC_20_in2_ready;
	wire branchC_20_in2_valid;
	wire [0 : 0]branchC_20_out1_data;
	wire branchC_20_out1_ready;
	wire branchC_20_out1_valid;
	wire [0 : 0]branchC_20_out2_data;
	wire branchC_20_out2_ready;
	wire branchC_20_out2_valid;

	wire fork_25_clk;
	wire fork_25_rst;
	wire [0 : 0]fork_25_in1_data;
	wire fork_25_in1_ready;
	wire fork_25_in1_valid;
	wire [0 : 0]fork_25_out1_data;
	wire fork_25_out1_ready;
	wire fork_25_out1_valid;
	wire [0 : 0]fork_25_out2_data;
	wire fork_25_out2_ready;
	wire fork_25_out2_valid;

	wire source_9_clk;
	wire source_9_rst;
	wire [0 : 0]source_9_out1_data;
	wire source_9_out1_ready;
	wire source_9_out1_valid;

	wire source_10_clk;
	wire source_10_rst;
	wire [4 : 0]source_10_out1_data;
	wire source_10_out1_ready;
	wire source_10_out1_valid;

	wire ret_0_clk;
	wire ret_0_rst;
	wire [0 : 0]ret_0_in1_data;
	wire ret_0_in1_ready;
	wire ret_0_in1_valid;
	wire [0 : 0]ret_0_out1_data;
	wire ret_0_out1_ready;
	wire ret_0_out1_valid;

	wire end_0_clk;
	wire end_0_rst;
	wire [0 : 0]end_0_in1_data;
	wire end_0_in1_ready;
	wire end_0_in1_valid;
	wire [0 : 0]end_0_in2_data;
	wire end_0_in2_ready;
	wire end_0_in2_valid;
	wire [0 : 0]end_0_in3_data;
	wire end_0_in3_ready;
	wire end_0_in3_valid;
	wire [0 : 0]end_0_out1_data;
	wire end_0_out1_ready;
	wire end_0_out1_valid;

	wire phiC_14_clk;
	wire phiC_14_rst;
	wire [0 : 0]phiC_14_in1_data;
	wire phiC_14_in1_ready;
	wire phiC_14_in1_valid;
	wire [0 : 0]phiC_14_out1_data;
	wire phiC_14_out1_ready;
	wire phiC_14_out1_valid;

	wire phi_6_clk;
	wire phi_6_rst;
	wire [0 : 0]phi_6_in1_data;
	wire phi_6_in1_ready;
	wire phi_6_in1_valid;
	wire [4 : 0]phi_6_in2_data;
	wire phi_6_in2_ready;
	wire phi_6_in2_valid;
	wire [4 : 0]phi_6_in3_data;
	wire phi_6_in3_ready;
	wire phi_6_in3_valid;
	wire [4 : 0]phi_6_out1_data;
	wire phi_6_out1_ready;
	wire phi_6_out1_valid;

	wire brCst_block4_clk;
	wire brCst_block4_rst;
	wire [0 : 0]brCst_block4_in1_data;
	wire brCst_block4_in1_ready;
	wire brCst_block4_in1_valid;
	wire [0 : 0]brCst_block4_out1_data;
	wire brCst_block4_out1_ready;
	wire brCst_block4_out1_valid;

	wire cst_3_clk;
	wire cst_3_rst;
	wire [0 : 0]cst_3_in1_data;
	wire cst_3_in1_ready;
	wire cst_3_in1_valid;
	wire [0 : 0]cst_3_out1_data;
	wire cst_3_out1_ready;
	wire cst_3_out1_valid;

	wire phi_n3_clk;
	wire phi_n3_rst;
	wire [4 : 0]phi_n3_in1_data;
	wire phi_n3_in1_ready;
	wire phi_n3_in1_valid;
	wire [4 : 0]phi_n3_in2_data;
	wire phi_n3_in2_ready;
	wire phi_n3_in2_valid;
	wire [4 : 0]phi_n3_out1_data;
	wire phi_n3_out1_ready;
	wire phi_n3_out1_valid;

	wire branch_5_clk;
	wire branch_5_rst;
	wire [0 : 0]branch_5_in1_data;
	wire branch_5_in1_ready;
	wire branch_5_in1_valid;
	wire [0 : 0]branch_5_in2_data;
	wire branch_5_in2_ready;
	wire branch_5_in2_valid;
	wire [0 : 0]branch_5_out1_data;
	wire branch_5_out1_ready;
	wire branch_5_out1_valid;
	wire [0 : 0]branch_5_out2_data;
	wire branch_5_out2_ready;
	wire branch_5_out2_valid;

	wire branch_6_clk;
	wire branch_6_rst;
	wire [4 : 0]branch_6_in1_data;
	wire branch_6_in1_ready;
	wire branch_6_in1_valid;
	wire [0 : 0]branch_6_in2_data;
	wire branch_6_in2_ready;
	wire branch_6_in2_valid;
	wire [4 : 0]branch_6_out1_data;
	wire branch_6_out1_ready;
	wire branch_6_out1_valid;
	wire [4 : 0]branch_6_out2_data;
	wire branch_6_out2_ready;
	wire branch_6_out2_valid;

	wire branch_7_clk;
	wire branch_7_rst;
	wire [4 : 0]branch_7_in1_data;
	wire branch_7_in1_ready;
	wire branch_7_in1_valid;
	wire [0 : 0]branch_7_in2_data;
	wire branch_7_in2_ready;
	wire branch_7_in2_valid;
	wire [4 : 0]branch_7_out1_data;
	wire branch_7_out1_ready;
	wire branch_7_out1_valid;
	wire [4 : 0]branch_7_out2_data;
	wire branch_7_out2_ready;
	wire branch_7_out2_valid;

	wire fork_12_clk;
	wire fork_12_rst;
	wire [0 : 0]fork_12_in1_data;
	wire fork_12_in1_ready;
	wire fork_12_in1_valid;
	wire [0 : 0]fork_12_out1_data;
	wire fork_12_out1_ready;
	wire fork_12_out1_valid;
	wire [0 : 0]fork_12_out2_data;
	wire fork_12_out2_ready;
	wire fork_12_out2_valid;
	wire [0 : 0]fork_12_out3_data;
	wire fork_12_out3_ready;
	wire fork_12_out3_valid;
	wire [0 : 0]fork_12_out4_data;
	wire fork_12_out4_ready;
	wire fork_12_out4_valid;

	wire phiC_10_clk;
	wire phiC_10_rst;
	wire [0 : 0]phiC_10_in1_data;
	wire phiC_10_in1_ready;
	wire phiC_10_in1_valid;
	wire [0 : 0]phiC_10_in2_data;
	wire phiC_10_in2_ready;
	wire phiC_10_in2_valid;
	wire [0 : 0]phiC_10_out1_data;
	wire phiC_10_out1_ready;
	wire phiC_10_out1_valid;
	wire [0 : 0]phiC_10_out2_data;
	wire phiC_10_out2_ready;
	wire phiC_10_out2_valid;

	wire forkC_21_clk;
	wire forkC_21_rst;
	wire [0 : 0]forkC_21_in1_data;
	wire forkC_21_in1_ready;
	wire forkC_21_in1_valid;
	wire [0 : 0]forkC_21_out1_data;
	wire forkC_21_out1_ready;
	wire forkC_21_out1_valid;
	wire [0 : 0]forkC_21_out2_data;
	wire forkC_21_out2_ready;
	wire forkC_21_out2_valid;
	wire [0 : 0]forkC_21_out3_data;
	wire forkC_21_out3_ready;
	wire forkC_21_out3_valid;

	wire branchC_17_clk;
	wire branchC_17_rst;
	wire [0 : 0]branchC_17_in1_data;
	wire branchC_17_in1_ready;
	wire branchC_17_in1_valid;
	wire [0 : 0]branchC_17_in2_data;
	wire branchC_17_in2_ready;
	wire branchC_17_in2_valid;
	wire [0 : 0]branchC_17_out1_data;
	wire branchC_17_out1_ready;
	wire branchC_17_out1_valid;
	wire [0 : 0]branchC_17_out2_data;
	wire branchC_17_out2_ready;
	wire branchC_17_out2_valid;

	wire phi_8_clk;
	wire phi_8_rst;
	wire [0 : 0]phi_8_in1_data;
	wire phi_8_in1_ready;
	wire phi_8_in1_valid;
	wire [4 : 0]phi_8_in2_data;
	wire phi_8_in2_ready;
	wire phi_8_in2_valid;
	wire [4 : 0]phi_8_in3_data;
	wire phi_8_in3_ready;
	wire phi_8_in3_valid;
	wire [4 : 0]phi_8_out1_data;
	wire phi_8_out1_ready;
	wire phi_8_out1_valid;

	wire cst_4_clk;
	wire cst_4_rst;
	wire [2 : 0]cst_4_in1_data;
	wire cst_4_in1_ready;
	wire cst_4_in1_valid;
	wire [2 : 0]cst_4_out1_data;
	wire cst_4_out1_ready;
	wire cst_4_out1_valid;

	wire shl_9_clk;
	wire shl_9_rst;
	wire [8 : 0]shl_9_in1_data;
	wire shl_9_in1_ready;
	wire shl_9_in1_valid;
	wire [8 : 0]shl_9_in2_data;
	wire shl_9_in2_ready;
	wire shl_9_in2_valid;
	wire [8 : 0]shl_9_out1_data;
	wire shl_9_out1_ready;
	wire shl_9_out1_valid;

	wire add_10_clk;
	wire add_10_rst;
	wire [9 : 0]add_10_in1_data;
	wire add_10_in1_ready;
	wire add_10_in1_valid;
	wire [9 : 0]add_10_in2_data;
	wire add_10_in2_ready;
	wire add_10_in2_valid;
	wire [9 : 0]add_10_out1_data;
	wire add_10_out1_ready;
	wire add_10_out1_valid;

	wire load_13_clk;
	wire load_13_rst;
	wire [31 : 0]load_13_in1_data;
	wire load_13_in1_ready;
	wire load_13_in1_valid;
	wire [9 : 0]load_13_in2_data;
	wire load_13_in2_ready;
	wire load_13_in2_valid;
	wire [31 : 0]load_13_out1_data;
	wire load_13_out1_ready;
	wire load_13_out1_valid;
	wire [9 : 0]load_13_out2_data;
	wire load_13_out2_ready;
	wire load_13_out2_valid;

	wire load_16_clk;
	wire load_16_rst;
	wire [31 : 0]load_16_in1_data;
	wire load_16_in1_ready;
	wire load_16_in1_valid;
	wire [4 : 0]load_16_in2_data;
	wire load_16_in2_ready;
	wire load_16_in2_valid;
	wire [31 : 0]load_16_out1_data;
	wire load_16_out1_ready;
	wire load_16_out1_valid;
	wire [4 : 0]load_16_out2_data;
	wire load_16_out2_ready;
	wire load_16_out2_valid;

	wire cst_5_clk;
	wire cst_5_rst;
	wire [2 : 0]cst_5_in1_data;
	wire cst_5_in1_ready;
	wire cst_5_in1_valid;
	wire [2 : 0]cst_5_out1_data;
	wire cst_5_out1_ready;
	wire cst_5_out1_valid;

	wire shl_17_clk;
	wire shl_17_rst;
	wire [8 : 0]shl_17_in1_data;
	wire shl_17_in1_ready;
	wire shl_17_in1_valid;
	wire [8 : 0]shl_17_in2_data;
	wire shl_17_in2_ready;
	wire shl_17_in2_valid;
	wire [8 : 0]shl_17_out1_data;
	wire shl_17_out1_ready;
	wire shl_17_out1_valid;

	wire add_18_clk;
	wire add_18_rst;
	wire [9 : 0]add_18_in1_data;
	wire add_18_in1_ready;
	wire add_18_in1_valid;
	wire [9 : 0]add_18_in2_data;
	wire add_18_in2_ready;
	wire add_18_in2_valid;
	wire [9 : 0]add_18_out1_data;
	wire add_18_out1_ready;
	wire add_18_out1_valid;

	wire load_21_clk;
	wire load_21_rst;
	wire [31 : 0]load_21_in1_data;
	wire load_21_in1_ready;
	wire load_21_in1_valid;
	wire [9 : 0]load_21_in2_data;
	wire load_21_in2_ready;
	wire load_21_in2_valid;
	wire [31 : 0]load_21_out1_data;
	wire load_21_out1_ready;
	wire load_21_out1_valid;
	wire [9 : 0]load_21_out2_data;
	wire load_21_out2_ready;
	wire load_21_out2_valid;

	wire mul_22_clk;
	wire mul_22_rst;
	wire [15 : 0]mul_22_in1_data;
	wire mul_22_in1_ready;
	wire mul_22_in1_valid;
	wire [15 : 0]mul_22_in2_data;
	wire mul_22_in2_ready;
	wire mul_22_in2_valid;
	wire [31 : 0]mul_22_out1_data;
	wire mul_22_out1_ready;
	wire mul_22_out1_valid;

	wire sub_23_clk;
	wire sub_23_rst;
	wire [31 : 0]sub_23_in1_data;
	wire sub_23_in1_ready;
	wire sub_23_in1_valid;
	wire [31 : 0]sub_23_in2_data;
	wire sub_23_in2_ready;
	wire sub_23_in2_valid;
	wire [31 : 0]sub_23_out1_data;
	wire sub_23_out1_ready;
	wire sub_23_out1_valid;

	wire cst_6_clk;
	wire cst_6_rst;
	wire [2 : 0]cst_6_in1_data;
	wire cst_6_in1_ready;
	wire cst_6_in1_valid;
	wire [2 : 0]cst_6_out1_data;
	wire cst_6_out1_ready;
	wire cst_6_out1_valid;

	wire shl_24_clk;
	wire shl_24_rst;
	wire [8 : 0]shl_24_in1_data;
	wire shl_24_in1_ready;
	wire shl_24_in1_valid;
	wire [8 : 0]shl_24_in2_data;
	wire shl_24_in2_ready;
	wire shl_24_in2_valid;
	wire [8 : 0]shl_24_out1_data;
	wire shl_24_out1_ready;
	wire shl_24_out1_valid;

	wire add_25_clk;
	wire add_25_rst;
	wire [9 : 0]add_25_in1_data;
	wire add_25_in1_ready;
	wire add_25_in1_valid;
	wire [9 : 0]add_25_in2_data;
	wire add_25_in2_ready;
	wire add_25_in2_valid;
	wire [9 : 0]add_25_out1_data;
	wire add_25_out1_ready;
	wire add_25_out1_valid;

	wire store_0_clk;
	wire store_0_rst;
	wire [31 : 0]store_0_in1_data;
	wire store_0_in1_ready;
	wire store_0_in1_valid;
	wire [9 : 0]store_0_in2_data;
	wire store_0_in2_ready;
	wire store_0_in2_valid;
	wire [31 : 0]store_0_out1_data;
	wire store_0_out1_ready;
	wire store_0_out1_valid;
	wire [9 : 0]store_0_out2_data;
	wire store_0_out2_ready;
	wire store_0_out2_valid;

	wire cst_7_clk;
	wire cst_7_rst;
	wire [0 : 0]cst_7_in1_data;
	wire cst_7_in1_ready;
	wire cst_7_in1_valid;
	wire [0 : 0]cst_7_out1_data;
	wire cst_7_out1_ready;
	wire cst_7_out1_valid;

	wire add_28_clk;
	wire add_28_rst;
	wire [4 : 0]add_28_in1_data;
	wire add_28_in1_ready;
	wire add_28_in1_valid;
	wire [4 : 0]add_28_in2_data;
	wire add_28_in2_ready;
	wire add_28_in2_valid;
	wire [4 : 0]add_28_out1_data;
	wire add_28_out1_ready;
	wire add_28_out1_valid;

	wire cst_8_clk;
	wire cst_8_rst;
	wire [4 : 0]cst_8_in1_data;
	wire cst_8_in1_ready;
	wire cst_8_in1_valid;
	wire [4 : 0]cst_8_out1_data;
	wire cst_8_out1_ready;
	wire cst_8_out1_valid;

	wire icmp_29_clk;
	wire icmp_29_rst;
	wire [4 : 0]icmp_29_in1_data;
	wire icmp_29_in1_ready;
	wire icmp_29_in1_valid;
	wire [4 : 0]icmp_29_in2_data;
	wire icmp_29_in2_ready;
	wire icmp_29_in2_valid;
	wire [0 : 0]icmp_29_out1_data;
	wire icmp_29_out1_ready;
	wire icmp_29_out1_valid;

	wire phi_n6_clk;
	wire phi_n6_rst;
	wire [4 : 0]phi_n6_in1_data;
	wire phi_n6_in1_ready;
	wire phi_n6_in1_valid;
	wire [4 : 0]phi_n6_in2_data;
	wire phi_n6_in2_ready;
	wire phi_n6_in2_valid;
	wire [4 : 0]phi_n6_out1_data;
	wire phi_n6_out1_ready;
	wire phi_n6_out1_valid;

	wire phi_n7_clk;
	wire phi_n7_rst;
	wire [4 : 0]phi_n7_in1_data;
	wire phi_n7_in1_ready;
	wire phi_n7_in1_valid;
	wire [4 : 0]phi_n7_in2_data;
	wire phi_n7_in2_ready;
	wire phi_n7_in2_valid;
	wire [4 : 0]phi_n7_out1_data;
	wire phi_n7_out1_ready;
	wire phi_n7_out1_valid;

	wire fork_2_clk;
	wire fork_2_rst;
	wire [4 : 0]fork_2_in1_data;
	wire fork_2_in1_ready;
	wire fork_2_in1_valid;
	wire [4 : 0]fork_2_out1_data;
	wire fork_2_out1_ready;
	wire fork_2_out1_valid;
	wire [4 : 0]fork_2_out2_data;
	wire fork_2_out2_ready;
	wire fork_2_out2_valid;
	wire [4 : 0]fork_2_out3_data;
	wire fork_2_out3_ready;
	wire fork_2_out3_valid;
	wire [4 : 0]fork_2_out4_data;
	wire fork_2_out4_ready;
	wire fork_2_out4_valid;

	wire fork_3_clk;
	wire fork_3_rst;
	wire [4 : 0]fork_3_in1_data;
	wire fork_3_in1_ready;
	wire fork_3_in1_valid;
	wire [4 : 0]fork_3_out1_data;
	wire fork_3_out1_ready;
	wire fork_3_out1_valid;
	wire [4 : 0]fork_3_out2_data;
	wire fork_3_out2_ready;
	wire fork_3_out2_valid;

	wire fork_7_clk;
	wire fork_7_rst;
	wire [4 : 0]fork_7_in1_data;
	wire fork_7_in1_ready;
	wire fork_7_in1_valid;
	wire [4 : 0]fork_7_out1_data;
	wire fork_7_out1_ready;
	wire fork_7_out1_valid;
	wire [4 : 0]fork_7_out2_data;
	wire fork_7_out2_ready;
	wire fork_7_out2_valid;
	wire [4 : 0]fork_7_out3_data;
	wire fork_7_out3_ready;
	wire fork_7_out3_valid;

	wire fork_8_clk;
	wire fork_8_rst;
	wire [4 : 0]fork_8_in1_data;
	wire fork_8_in1_ready;
	wire fork_8_in1_valid;
	wire [4 : 0]fork_8_out1_data;
	wire fork_8_out1_ready;
	wire fork_8_out1_valid;
	wire [4 : 0]fork_8_out2_data;
	wire fork_8_out2_ready;
	wire fork_8_out2_valid;
	wire [4 : 0]fork_8_out3_data;
	wire fork_8_out3_ready;
	wire fork_8_out3_valid;

	wire branch_8_clk;
	wire branch_8_rst;
	wire [4 : 0]branch_8_in1_data;
	wire branch_8_in1_ready;
	wire branch_8_in1_valid;
	wire [0 : 0]branch_8_in2_data;
	wire branch_8_in2_ready;
	wire branch_8_in2_valid;
	wire [4 : 0]branch_8_out1_data;
	wire branch_8_out1_ready;
	wire branch_8_out1_valid;
	wire [4 : 0]branch_8_out2_data;
	wire branch_8_out2_ready;
	wire branch_8_out2_valid;

	wire branch_9_clk;
	wire branch_9_rst;
	wire [4 : 0]branch_9_in1_data;
	wire branch_9_in1_ready;
	wire branch_9_in1_valid;
	wire [0 : 0]branch_9_in2_data;
	wire branch_9_in2_ready;
	wire branch_9_in2_valid;
	wire [4 : 0]branch_9_out1_data;
	wire branch_9_out1_ready;
	wire branch_9_out1_valid;
	wire [4 : 0]branch_9_out2_data;
	wire branch_9_out2_ready;
	wire branch_9_out2_valid;

	wire branch_10_clk;
	wire branch_10_rst;
	wire [4 : 0]branch_10_in1_data;
	wire branch_10_in1_ready;
	wire branch_10_in1_valid;
	wire [0 : 0]branch_10_in2_data;
	wire branch_10_in2_ready;
	wire branch_10_in2_valid;
	wire [4 : 0]branch_10_out1_data;
	wire branch_10_out1_ready;
	wire branch_10_out1_valid;
	wire [4 : 0]branch_10_out2_data;
	wire branch_10_out2_ready;
	wire branch_10_out2_valid;

	wire fork_13_clk;
	wire fork_13_rst;
	wire [0 : 0]fork_13_in1_data;
	wire fork_13_in1_ready;
	wire fork_13_in1_valid;
	wire [0 : 0]fork_13_out1_data;
	wire fork_13_out1_ready;
	wire fork_13_out1_valid;
	wire [0 : 0]fork_13_out2_data;
	wire fork_13_out2_ready;
	wire fork_13_out2_valid;
	wire [0 : 0]fork_13_out3_data;
	wire fork_13_out3_ready;
	wire fork_13_out3_valid;
	wire [0 : 0]fork_13_out4_data;
	wire fork_13_out4_ready;
	wire fork_13_out4_valid;

	wire cst_13_clk;
	wire cst_13_rst;
	wire [0 : 0]cst_13_in1_data;
	wire cst_13_in1_ready;
	wire cst_13_in1_valid;
	wire [0 : 0]cst_13_out1_data;
	wire cst_13_out1_ready;
	wire cst_13_out1_valid;

	wire phiC_11_clk;
	wire phiC_11_rst;
	wire [0 : 0]phiC_11_in1_data;
	wire phiC_11_in1_ready;
	wire phiC_11_in1_valid;
	wire [0 : 0]phiC_11_in2_data;
	wire phiC_11_in2_ready;
	wire phiC_11_in2_valid;
	wire [0 : 0]phiC_11_out1_data;
	wire phiC_11_out1_ready;
	wire phiC_11_out1_valid;
	wire [0 : 0]phiC_11_out2_data;
	wire phiC_11_out2_ready;
	wire phiC_11_out2_valid;

	wire forkC_22_clk;
	wire forkC_22_rst;
	wire [0 : 0]forkC_22_in1_data;
	wire forkC_22_in1_ready;
	wire forkC_22_in1_valid;
	wire [0 : 0]forkC_22_out1_data;
	wire forkC_22_out1_ready;
	wire forkC_22_out1_valid;
	wire [0 : 0]forkC_22_out2_data;
	wire forkC_22_out2_ready;
	wire forkC_22_out2_valid;

	wire branchC_18_clk;
	wire branchC_18_rst;
	wire [0 : 0]branchC_18_in1_data;
	wire branchC_18_in1_ready;
	wire branchC_18_in1_valid;
	wire [0 : 0]branchC_18_in2_data;
	wire branchC_18_in2_ready;
	wire branchC_18_in2_valid;
	wire [0 : 0]branchC_18_out1_data;
	wire branchC_18_out1_ready;
	wire branchC_18_out1_valid;
	wire [0 : 0]branchC_18_out2_data;
	wire branchC_18_out2_ready;
	wire branchC_18_out2_valid;

	wire source_2_clk;
	wire source_2_rst;
	wire [2 : 0]source_2_out1_data;
	wire source_2_out1_ready;
	wire source_2_out1_valid;

	wire source_3_clk;
	wire source_3_rst;
	wire [2 : 0]source_3_out1_data;
	wire source_3_out1_ready;
	wire source_3_out1_valid;

	wire source_4_clk;
	wire source_4_rst;
	wire [2 : 0]source_4_out1_data;
	wire source_4_out1_ready;
	wire source_4_out1_valid;

	wire source_5_clk;
	wire source_5_rst;
	wire [0 : 0]source_5_out1_data;
	wire source_5_out1_ready;
	wire source_5_out1_valid;

	wire source_6_clk;
	wire source_6_rst;
	wire [4 : 0]source_6_out1_data;
	wire source_6_out1_ready;
	wire source_6_out1_valid;

	wire phi_1_clk;
	wire phi_1_rst;
	wire [0 : 0]phi_1_in1_data;
	wire phi_1_in1_ready;
	wire phi_1_in1_valid;
	wire [4 : 0]phi_1_in2_data;
	wire phi_1_in2_ready;
	wire phi_1_in2_valid;
	wire [4 : 0]phi_1_in3_data;
	wire phi_1_in3_ready;
	wire phi_1_in3_valid;
	wire [4 : 0]phi_1_out1_data;
	wire phi_1_out1_ready;
	wire phi_1_out1_valid;

	wire cst_1_clk;
	wire cst_1_rst;
	wire [0 : 0]cst_1_in1_data;
	wire cst_1_in1_ready;
	wire cst_1_in1_valid;
	wire [0 : 0]cst_1_out1_data;
	wire cst_1_out1_ready;
	wire cst_1_out1_valid;

	wire add_2_clk;
	wire add_2_rst;
	wire [5 : 0]add_2_in1_data;
	wire add_2_in1_ready;
	wire add_2_in1_valid;
	wire [5 : 0]add_2_in2_data;
	wire add_2_in2_ready;
	wire add_2_in2_valid;
	wire [5 : 0]add_2_out1_data;
	wire add_2_out1_ready;
	wire add_2_out1_valid;

	wire cst_2_clk;
	wire cst_2_rst;
	wire [4 : 0]cst_2_in1_data;
	wire cst_2_in1_ready;
	wire cst_2_in1_valid;
	wire [4 : 0]cst_2_out1_data;
	wire cst_2_out1_ready;
	wire cst_2_out1_valid;

	wire icmp_3_clk;
	wire icmp_3_rst;
	wire [5 : 0]icmp_3_in1_data;
	wire icmp_3_in1_ready;
	wire icmp_3_in1_valid;
	wire [5 : 0]icmp_3_in2_data;
	wire icmp_3_in2_ready;
	wire icmp_3_in2_valid;
	wire [0 : 0]icmp_3_out1_data;
	wire icmp_3_out1_ready;
	wire icmp_3_out1_valid;

	wire fork_0_clk;
	wire fork_0_rst;
	wire [4 : 0]fork_0_in1_data;
	wire fork_0_in1_ready;
	wire fork_0_in1_valid;
	wire [4 : 0]fork_0_out1_data;
	wire fork_0_out1_ready;
	wire fork_0_out1_valid;
	wire [4 : 0]fork_0_out2_data;
	wire fork_0_out2_ready;
	wire fork_0_out2_valid;

	wire fork_1_clk;
	wire fork_1_rst;
	wire [5 : 0]fork_1_in1_data;
	wire fork_1_in1_ready;
	wire fork_1_in1_valid;
	wire [5 : 0]fork_1_out1_data;
	wire fork_1_out1_ready;
	wire fork_1_out1_valid;
	wire [5 : 0]fork_1_out2_data;
	wire fork_1_out2_ready;
	wire fork_1_out2_valid;

	wire branch_1_clk;
	wire branch_1_rst;
	wire [4 : 0]branch_1_in1_data;
	wire branch_1_in1_ready;
	wire branch_1_in1_valid;
	wire [0 : 0]branch_1_in2_data;
	wire branch_1_in2_ready;
	wire branch_1_in2_valid;
	wire [4 : 0]branch_1_out1_data;
	wire branch_1_out1_ready;
	wire branch_1_out1_valid;
	wire [4 : 0]branch_1_out2_data;
	wire branch_1_out2_ready;
	wire branch_1_out2_valid;

	wire branch_2_clk;
	wire branch_2_rst;
	wire [5 : 0]branch_2_in1_data;
	wire branch_2_in1_ready;
	wire branch_2_in1_valid;
	wire [0 : 0]branch_2_in2_data;
	wire branch_2_in2_ready;
	wire branch_2_in2_valid;
	wire [5 : 0]branch_2_out1_data;
	wire branch_2_out1_ready;
	wire branch_2_out1_valid;
	wire [5 : 0]branch_2_out2_data;
	wire branch_2_out2_ready;
	wire branch_2_out2_valid;

	wire fork_10_clk;
	wire fork_10_rst;
	wire [0 : 0]fork_10_in1_data;
	wire fork_10_in1_ready;
	wire fork_10_in1_valid;
	wire [0 : 0]fork_10_out1_data;
	wire fork_10_out1_ready;
	wire fork_10_out1_valid;
	wire [0 : 0]fork_10_out2_data;
	wire fork_10_out2_ready;
	wire fork_10_out2_valid;
	wire [0 : 0]fork_10_out3_data;
	wire fork_10_out3_ready;
	wire fork_10_out3_valid;

	wire phiC_8_clk;
	wire phiC_8_rst;
	wire [0 : 0]phiC_8_in1_data;
	wire phiC_8_in1_ready;
	wire phiC_8_in1_valid;
	wire [0 : 0]phiC_8_in2_data;
	wire phiC_8_in2_ready;
	wire phiC_8_in2_valid;
	wire [0 : 0]phiC_8_out1_data;
	wire phiC_8_out1_ready;
	wire phiC_8_out1_valid;
	wire [0 : 0]phiC_8_out2_data;
	wire phiC_8_out2_ready;
	wire phiC_8_out2_valid;

	wire branchC_15_clk;
	wire branchC_15_rst;
	wire [0 : 0]branchC_15_in1_data;
	wire branchC_15_in1_ready;
	wire branchC_15_in1_valid;
	wire [0 : 0]branchC_15_in2_data;
	wire branchC_15_in2_ready;
	wire branchC_15_in2_valid;
	wire [0 : 0]branchC_15_out1_data;
	wire branchC_15_out1_ready;
	wire branchC_15_out1_valid;
	wire [0 : 0]branchC_15_out2_data;
	wire branchC_15_out2_ready;
	wire branchC_15_out2_valid;

	wire source_0_clk;
	wire source_0_rst;
	wire [0 : 0]source_0_out1_data;
	wire source_0_out1_ready;
	wire source_0_out1_valid;

	wire source_1_clk;
	wire source_1_rst;
	wire [4 : 0]source_1_out1_data;
	wire source_1_out1_ready;
	wire source_1_out1_valid;

	wire MC_A_clk;
	wire MC_A_rst;
	wire [31 : 0]MC_A_in1_data;
	wire MC_A_in1_ready;
	wire MC_A_in1_valid;
	wire [9 : 0]MC_A_in2_data;
	wire MC_A_in2_ready;
	wire MC_A_in2_valid;
	wire [9 : 0]MC_A_in3_data;
	wire MC_A_in3_ready;
	wire MC_A_in3_valid;
	wire [9 : 0]MC_A_in4_data;
	wire MC_A_in4_ready;
	wire MC_A_in4_valid;
	wire [31 : 0]MC_A_in5_data;
	wire MC_A_in5_ready;
	wire MC_A_in5_valid;
	wire [31 : 0]MC_A_out1_data;
	wire MC_A_out1_ready;
	wire MC_A_out1_valid;
	wire [31 : 0]MC_A_out2_data;
	wire MC_A_out2_ready;
	wire MC_A_out2_valid;
	wire [0 : 0]MC_A_out3_data;
	wire MC_A_out3_ready;
	wire MC_A_out3_valid;

	wire MC_c_clk;
	wire MC_c_rst;
	wire [4 : 0]MC_c_in1_data;
	wire MC_c_in1_ready;
	wire MC_c_in1_valid;
	wire [31 : 0]MC_c_in2_data;
	wire MC_c_in2_ready;
	wire MC_c_in2_valid;
	wire [4 : 0]MC_c_in3_data;
	wire MC_c_in3_ready;
	wire MC_c_in3_valid;
	wire [31 : 0]MC_c_in4_data;
	wire MC_c_in4_ready;
	wire MC_c_in4_valid;
	wire [31 : 0]MC_c_out1_data;
	wire MC_c_out1_ready;
	wire MC_c_out1_valid;
	wire [0 : 0]MC_c_out2_data;
	wire MC_c_out2_ready;
	wire MC_c_out2_valid;

	wire sink_0_clk;
	wire sink_0_rst;
	wire [0 : 0]sink_0_in1_data;
	wire sink_0_in1_ready;
	wire sink_0_in1_valid;

	wire sink_1_clk;
	wire sink_1_rst;
	wire [5 : 0]sink_1_in1_data;
	wire sink_1_in1_ready;
	wire sink_1_in1_valid;

	wire sink_2_clk;
	wire sink_2_rst;
	wire [5 : 0]sink_2_in1_data;
	wire sink_2_in1_ready;
	wire sink_2_in1_valid;

	wire sink_3_clk;
	wire sink_3_rst;
	wire [4 : 0]sink_3_in1_data;
	wire sink_3_in1_ready;
	wire sink_3_in1_valid;

	wire sink_4_clk;
	wire sink_4_rst;
	wire [0 : 0]sink_4_in1_data;
	wire sink_4_in1_ready;
	wire sink_4_in1_valid;

	wire sink_5_clk;
	wire sink_5_rst;
	wire [4 : 0]sink_5_in1_data;
	wire sink_5_in1_ready;
	wire sink_5_in1_valid;

	wire sink_6_clk;
	wire sink_6_rst;
	wire [4 : 0]sink_6_in1_data;
	wire sink_6_in1_ready;
	wire sink_6_in1_valid;

	wire sink_7_clk;
	wire sink_7_rst;
	wire [4 : 0]sink_7_in1_data;
	wire sink_7_in1_ready;
	wire sink_7_in1_valid;

	wire sink_8_clk;
	wire sink_8_rst;
	wire [4 : 0]sink_8_in1_data;
	wire sink_8_in1_ready;
	wire sink_8_in1_valid;

	wire sink_9_clk;
	wire sink_9_rst;
	wire [4 : 0]sink_9_in1_data;
	wire sink_9_in1_ready;
	wire sink_9_in1_valid;

	wire sink_10_clk;
	wire sink_10_rst;
	wire [0 : 0]sink_10_in1_data;
	wire sink_10_in1_ready;
	wire sink_10_in1_valid;

	wire sink_11_clk;
	wire sink_11_rst;
	wire [0 : 0]sink_11_in1_data;
	wire sink_11_in1_ready;
	wire sink_11_in1_valid;

	wire sink_12_clk;
	wire sink_12_rst;
	wire [0 : 0]sink_12_in1_data;
	wire sink_12_in1_ready;
	wire sink_12_in1_valid;

	wire Buffer_100_clk;
	wire Buffer_100_rst;
	wire [31 : 0]Buffer_100_in1_data;
	wire Buffer_100_in1_ready;
	wire Buffer_100_in1_valid;
	wire [31 : 0]Buffer_100_out1_data;
	wire Buffer_100_out1_ready;
	wire Buffer_100_out1_valid;

	wire Buffer_101_clk;
	wire Buffer_101_rst;
	wire [31 : 0]Buffer_101_in1_data;
	wire Buffer_101_in1_ready;
	wire Buffer_101_in1_valid;
	wire [31 : 0]Buffer_101_out1_data;
	wire Buffer_101_out1_ready;
	wire Buffer_101_out1_valid;

	wire Buffer_102_clk;
	wire Buffer_102_rst;
	wire [31 : 0]Buffer_102_in1_data;
	wire Buffer_102_in1_ready;
	wire Buffer_102_in1_valid;
	wire [31 : 0]Buffer_102_out1_data;
	wire Buffer_102_out1_ready;
	wire Buffer_102_out1_valid;

	wire Buffer_103_clk;
	wire Buffer_103_rst;
	wire [31 : 0]Buffer_103_in1_data;
	wire Buffer_103_in1_ready;
	wire Buffer_103_in1_valid;
	wire [31 : 0]Buffer_103_out1_data;
	wire Buffer_103_out1_ready;
	wire Buffer_103_out1_valid;

	wire Buffer_104_clk;
	wire Buffer_104_rst;
	wire [31 : 0]Buffer_104_in1_data;
	wire Buffer_104_in1_ready;
	wire Buffer_104_in1_valid;
	wire [31 : 0]Buffer_104_out1_data;
	wire Buffer_104_out1_ready;
	wire Buffer_104_out1_valid;

	wire Buffer_105_clk;
	wire Buffer_105_rst;
	wire [31 : 0]Buffer_105_in1_data;
	wire Buffer_105_in1_ready;
	wire Buffer_105_in1_valid;
	wire [31 : 0]Buffer_105_out1_data;
	wire Buffer_105_out1_ready;
	wire Buffer_105_out1_valid;

	wire Buffer_106_clk;
	wire Buffer_106_rst;
	wire [31 : 0]Buffer_106_in1_data;
	wire Buffer_106_in1_ready;
	wire Buffer_106_in1_valid;
	wire [31 : 0]Buffer_106_out1_data;
	wire Buffer_106_out1_ready;
	wire Buffer_106_out1_valid;

	wire Buffer_107_clk;
	wire Buffer_107_rst;
	wire [31 : 0]Buffer_107_in1_data;
	wire Buffer_107_in1_ready;
	wire Buffer_107_in1_valid;
	wire [31 : 0]Buffer_107_out1_data;
	wire Buffer_107_out1_ready;
	wire Buffer_107_out1_valid;

	wire Buffer_108_clk;
	wire Buffer_108_rst;
	wire [31 : 0]Buffer_108_in1_data;
	wire Buffer_108_in1_ready;
	wire Buffer_108_in1_valid;
	wire [31 : 0]Buffer_108_out1_data;
	wire Buffer_108_out1_ready;
	wire Buffer_108_out1_valid;



	assign brCst_block1_clk = clk;
	assign brCst_block1_rst = rst;
	assign fork_18_in1_data = brCst_block1_out1_data;
	assign fork_18_in1_valid = brCst_block1_out1_valid;
	assign brCst_block1_out1_ready = fork_18_in1_ready;

	assign cst_0_clk = clk;
	assign cst_0_rst = rst;
	assign branch_0_in1_data = cst_0_out1_data;
	assign branch_0_in1_valid = cst_0_out1_valid;
	assign cst_0_out1_ready = branch_0_in1_ready;

	assign branch_0_clk = clk;
	assign branch_0_rst = rst;
	assign phi_1_in2_data = branch_0_out1_data;
	assign phi_1_in2_valid = branch_0_out1_valid;
	assign branch_0_out1_ready = phi_1_in2_ready;
	assign sink_0_in1_data = branch_0_out2_data;
	assign sink_0_in1_valid = branch_0_out2_valid;
	assign branch_0_out2_ready = sink_0_in1_ready;

	assign start_0_clk = clk;
	assign start_0_rst = rst;
	assign start_0_in1_data = start_in;
	assign start_0_in1_valid = start_valid;
	assign start_ready = start_0_in1_ready;
	assign forkC_17_in1_data = start_0_out1_data;
	assign forkC_17_in1_valid = start_0_out1_valid;
	assign start_0_out1_ready = forkC_17_in1_ready;

	assign forkC_17_clk = clk;
	assign forkC_17_rst = rst;
	assign cst_0_in1_data = forkC_17_out1_data;
	assign cst_0_in1_valid = forkC_17_out1_valid;
	assign forkC_17_out1_ready = cst_0_in1_ready;
	assign branchC_14_in1_data = forkC_17_out2_data;
	assign branchC_14_in1_valid = forkC_17_out2_valid;
	assign forkC_17_out2_ready = branchC_14_in1_ready;
	assign brCst_block1_in1_data = forkC_17_out3_data;
	assign brCst_block1_in1_valid = forkC_17_out3_valid;
	assign forkC_17_out3_ready = brCst_block1_in1_ready;

	assign branchC_14_clk = clk;
	assign branchC_14_rst = rst;
	assign phiC_8_in1_data = branchC_14_out1_data;
	assign phiC_8_in1_valid = branchC_14_out1_valid;
	assign branchC_14_out1_ready = phiC_8_in1_ready;
	assign sink_10_in1_data = branchC_14_out2_data;
	assign sink_10_in1_valid = branchC_14_out2_valid;
	assign branchC_14_out2_ready = sink_10_in1_ready;

	assign fork_18_clk = clk;
	assign fork_18_rst = rst;
	assign branch_0_in2_data = fork_18_out1_data;
	assign branch_0_in2_valid = fork_18_out1_valid;
	assign fork_18_out1_ready = branch_0_in2_ready;
	assign branchC_14_in2_data = fork_18_out2_data;
	assign branchC_14_in2_valid = fork_18_out2_valid;
	assign fork_18_out2_ready = branchC_14_in2_ready;

	assign brCst_block3_clk = clk;
	assign brCst_block3_rst = rst;
	assign fork_11_in1_data = brCst_block3_out1_data;
	assign fork_11_in1_valid = brCst_block3_out1_valid;
	assign brCst_block3_out1_ready = fork_11_in1_ready;

	assign phi_n1_clk = clk;
	assign phi_n1_rst = rst;
	assign branch_3_in1_data = phi_n1_out1_data;
	assign branch_3_in1_valid = phi_n1_out1_valid;
	assign phi_n1_out1_ready = branch_3_in1_ready;

	assign phi_n2_clk = clk;
	assign phi_n2_rst = rst;
	assign branch_4_in1_data = phi_n2_out1_data;
	assign branch_4_in1_valid = phi_n2_out1_valid;
	assign phi_n2_out1_ready = branch_4_in1_ready;

	assign branch_3_clk = clk;
	assign branch_3_rst = rst;
	assign phi_6_in2_data = branch_3_out1_data;
	assign phi_6_in2_valid = branch_3_out1_valid;
	assign branch_3_out1_ready = phi_6_in2_ready;
	assign sink_2_in1_data = branch_3_out2_data;
	assign sink_2_in1_valid = branch_3_out2_valid;
	assign branch_3_out2_ready = sink_2_in1_ready;

	assign branch_4_clk = clk;
	assign branch_4_rst = rst;
	assign phi_n3_in1_data = branch_4_out1_data;
	assign phi_n3_in1_valid = branch_4_out1_valid;
	assign branch_4_out1_ready = phi_n3_in1_ready;
	assign sink_3_in1_data = branch_4_out2_data;
	assign sink_3_in1_valid = branch_4_out2_valid;
	assign branch_4_out2_ready = sink_3_in1_ready;

	assign fork_11_clk = clk;
	assign fork_11_rst = rst;
	assign branch_4_in2_data = fork_11_out1_data;
	assign branch_4_in2_valid = fork_11_out1_valid;
	assign fork_11_out1_ready = branch_4_in2_ready;
	assign branch_3_in2_data = fork_11_out2_data;
	assign branch_3_in2_valid = fork_11_out2_valid;
	assign fork_11_out2_ready = branch_3_in2_ready;
	assign branchC_16_in2_data = fork_11_out3_data;
	assign branchC_16_in2_valid = fork_11_out3_valid;
	assign fork_11_out3_ready = branchC_16_in2_ready;

	assign phiC_9_clk = clk;
	assign phiC_9_rst = rst;
	assign forkC_20_in1_data = phiC_9_out1_data;
	assign forkC_20_in1_valid = phiC_9_out1_valid;
	assign phiC_9_out1_ready = forkC_20_in1_ready;

	assign forkC_20_clk = clk;
	assign forkC_20_rst = rst;
	assign branchC_16_in1_data = forkC_20_out1_data;
	assign branchC_16_in1_valid = forkC_20_out1_valid;
	assign forkC_20_out1_ready = branchC_16_in1_ready;
	assign brCst_block3_in1_data = forkC_20_out2_data;
	assign brCst_block3_in1_valid = forkC_20_out2_valid;
	assign forkC_20_out2_ready = brCst_block3_in1_ready;

	assign branchC_16_clk = clk;
	assign branchC_16_rst = rst;
	assign phiC_10_in1_data = branchC_16_out1_data;
	assign phiC_10_in1_valid = branchC_16_out1_valid;
	assign branchC_16_out1_ready = phiC_10_in1_ready;
	assign sink_11_in1_data = branchC_16_out2_data;
	assign sink_11_in1_valid = branchC_16_out2_valid;
	assign branchC_16_out2_ready = sink_11_in1_ready;

	assign cst_9_clk = clk;
	assign cst_9_rst = rst;
	assign add_31_in2_data = cst_9_out1_data;
	assign add_31_in2_valid = cst_9_out1_valid;
	assign cst_9_out1_ready = add_31_in2_ready;

	assign add_31_clk = clk;
	assign add_31_rst = rst;
	assign branch_11_in1_data = add_31_out1_data;
	assign branch_11_in1_valid = add_31_out1_valid;
	assign add_31_out1_ready = branch_11_in1_ready;

	assign cst_10_clk = clk;
	assign cst_10_rst = rst;
	assign icmp_32_in2_data = cst_10_out1_data;
	assign icmp_32_in2_valid = cst_10_out1_valid;
	assign cst_10_out1_ready = icmp_32_in2_ready;

	assign icmp_32_clk = clk;
	assign icmp_32_rst = rst;
	assign fork_14_in1_data = icmp_32_out1_data;
	assign fork_14_in1_valid = icmp_32_out1_valid;
	assign icmp_32_out1_ready = fork_14_in1_ready;

	assign phi_n4_clk = clk;
	assign phi_n4_rst = rst;
	assign fork_5_in1_data = phi_n4_out1_data;
	assign fork_5_in1_valid = phi_n4_out1_valid;
	assign phi_n4_out1_ready = fork_5_in1_ready;

	assign phi_n5_clk = clk;
	assign phi_n5_rst = rst;
	assign branch_12_in1_data = phi_n5_out1_data;
	assign branch_12_in1_valid = phi_n5_out1_valid;
	assign phi_n5_out1_ready = branch_12_in1_ready;

	assign fork_5_clk = clk;
	assign fork_5_rst = rst;
	assign add_31_in1_data = fork_5_out1_data;
	assign add_31_in1_valid = fork_5_out1_valid;
	assign fork_5_out1_ready = add_31_in1_ready;
	assign icmp_32_in1_data = fork_5_out2_data;
	assign icmp_32_in1_valid = fork_5_out2_valid;
	assign fork_5_out2_ready = icmp_32_in1_ready;

	assign branch_11_clk = clk;
	assign branch_11_rst = rst;
	assign Buffer_104_in1_data = branch_11_out1_data;
	assign Buffer_104_in1_valid = branch_11_out1_valid;
	assign branch_11_out1_ready = Buffer_104_in1_ready;
	assign sink_8_in1_data = branch_11_out2_data;
	assign sink_8_in1_valid = branch_11_out2_valid;
	assign branch_11_out2_ready = sink_8_in1_ready;

	assign branch_12_clk = clk;
	assign branch_12_rst = rst;
	assign Buffer_105_in1_data = branch_12_out1_data;
	assign Buffer_105_in1_valid = branch_12_out1_valid;
	assign branch_12_out1_ready = Buffer_105_in1_ready;
	assign phi_n0_in2_data = branch_12_out2_data;
	assign phi_n0_in2_valid = branch_12_out2_valid;
	assign branch_12_out2_ready = phi_n0_in2_ready;

	assign fork_14_clk = clk;
	assign fork_14_rst = rst;
	assign branch_12_in2_data = fork_14_out1_data;
	assign branch_12_in2_valid = fork_14_out1_valid;
	assign fork_14_out1_ready = branch_12_in2_ready;
	assign branch_11_in2_data = fork_14_out2_data;
	assign branch_11_in2_valid = fork_14_out2_valid;
	assign fork_14_out2_ready = branch_11_in2_ready;
	assign branchC_19_in2_data = fork_14_out3_data;
	assign branchC_19_in2_valid = fork_14_out3_valid;
	assign fork_14_out3_ready = branchC_19_in2_ready;

	assign phiC_12_clk = clk;
	assign phiC_12_rst = rst;
	assign branchC_19_in1_data = phiC_12_out1_data;
	assign branchC_19_in1_valid = phiC_12_out1_valid;
	assign phiC_12_out1_ready = branchC_19_in1_ready;

	assign branchC_19_clk = clk;
	assign branchC_19_rst = rst;
	assign Buffer_106_in1_data = branchC_19_out1_data;
	assign Buffer_106_in1_valid = branchC_19_out1_valid;
	assign branchC_19_out1_ready = Buffer_106_in1_ready;
	assign phiC_13_in2_data = branchC_19_out2_data;
	assign phiC_13_in2_valid = branchC_19_out2_valid;
	assign branchC_19_out2_ready = phiC_13_in2_ready;

	assign source_7_clk = clk;
	assign source_7_rst = rst;
	assign cst_9_in1_data = source_7_out1_data;
	assign cst_9_in1_valid = source_7_out1_valid;
	assign source_7_out1_ready = cst_9_in1_ready;

	assign source_8_clk = clk;
	assign source_8_rst = rst;
	assign cst_10_in1_data = source_8_out1_data;
	assign cst_10_in1_valid = source_8_out1_valid;
	assign source_8_out1_ready = cst_10_in1_ready;

	assign cst_11_clk = clk;
	assign cst_11_rst = rst;
	assign add_34_in2_data = cst_11_out1_data;
	assign add_34_in2_valid = cst_11_out1_valid;
	assign cst_11_out1_ready = add_34_in2_ready;

	assign add_34_clk = clk;
	assign add_34_rst = rst;
	assign fork_4_in1_data = add_34_out1_data;
	assign fork_4_in1_valid = add_34_out1_valid;
	assign add_34_out1_ready = fork_4_in1_ready;

	assign cst_12_clk = clk;
	assign cst_12_rst = rst;
	assign icmp_35_in2_data = cst_12_out1_data;
	assign icmp_35_in2_valid = cst_12_out1_valid;
	assign cst_12_out1_ready = icmp_35_in2_ready;

	assign icmp_35_clk = clk;
	assign icmp_35_rst = rst;
	assign fork_25_in1_data = icmp_35_out1_data;
	assign fork_25_in1_valid = icmp_35_out1_valid;
	assign icmp_35_out1_ready = fork_25_in1_ready;

	assign phi_n0_clk = clk;
	assign phi_n0_rst = rst;
	assign add_34_in1_data = phi_n0_out1_data;
	assign add_34_in1_valid = phi_n0_out1_valid;
	assign phi_n0_out1_ready = add_34_in1_ready;

	assign fork_4_clk = clk;
	assign fork_4_rst = rst;
	assign icmp_35_in1_data = fork_4_out1_data;
	assign icmp_35_in1_valid = fork_4_out1_valid;
	assign fork_4_out1_ready = icmp_35_in1_ready;
	assign branch_13_in1_data = fork_4_out2_data;
	assign branch_13_in1_valid = fork_4_out2_valid;
	assign fork_4_out2_ready = branch_13_in1_ready;

	assign branch_13_clk = clk;
	assign branch_13_rst = rst;
	assign Buffer_107_in1_data = branch_13_out1_data;
	assign Buffer_107_in1_valid = branch_13_out1_valid;
	assign branch_13_out1_ready = Buffer_107_in1_ready;
	assign sink_9_in1_data = branch_13_out2_data;
	assign sink_9_in1_valid = branch_13_out2_valid;
	assign branch_13_out2_ready = sink_9_in1_ready;

	assign phiC_13_clk = clk;
	assign phiC_13_rst = rst;
	assign branchC_20_in1_data = phiC_13_out1_data;
	assign branchC_20_in1_valid = phiC_13_out1_valid;
	assign phiC_13_out1_ready = branchC_20_in1_ready;

	assign branchC_20_clk = clk;
	assign branchC_20_rst = rst;
	assign Buffer_108_in1_data = branchC_20_out1_data;
	assign Buffer_108_in1_valid = branchC_20_out1_valid;
	assign branchC_20_out1_ready = Buffer_108_in1_ready;
	assign phiC_14_in1_data = branchC_20_out2_data;
	assign phiC_14_in1_valid = branchC_20_out2_valid;
	assign branchC_20_out2_ready = phiC_14_in1_ready;

	assign fork_25_clk = clk;
	assign fork_25_rst = rst;
	assign branch_13_in2_data = fork_25_out1_data;
	assign branch_13_in2_valid = fork_25_out1_valid;
	assign fork_25_out1_ready = branch_13_in2_ready;
	assign branchC_20_in2_data = fork_25_out2_data;
	assign branchC_20_in2_valid = fork_25_out2_valid;
	assign fork_25_out2_ready = branchC_20_in2_ready;

	assign source_9_clk = clk;
	assign source_9_rst = rst;
	assign cst_11_in1_data = source_9_out1_data;
	assign cst_11_in1_valid = source_9_out1_valid;
	assign source_9_out1_ready = cst_11_in1_ready;

	assign source_10_clk = clk;
	assign source_10_rst = rst;
	assign cst_12_in1_data = source_10_out1_data;
	assign cst_12_in1_valid = source_10_out1_valid;
	assign source_10_out1_ready = cst_12_in1_ready;

	assign ret_0_clk = clk;
	assign ret_0_rst = rst;
	assign end_0_in3_data = ret_0_out1_data;
	assign end_0_in3_valid = ret_0_out1_valid;
	assign ret_0_out1_ready = end_0_in3_ready;

	assign end_0_clk = clk;
	assign end_0_rst = rst;
	assign end_out = end_0_out1_data;
	assign end_0_out1_ready = end_ready;
	assign end_valid = end_0_out1_valid;

	assign phiC_14_clk = clk;
	assign phiC_14_rst = rst;
	assign ret_0_in1_data = phiC_14_out1_data;
	assign ret_0_in1_valid = phiC_14_out1_valid;
	assign phiC_14_out1_ready = ret_0_in1_ready;

	assign phi_6_clk = clk;
	assign phi_6_rst = rst;
	assign branch_6_in1_data = phi_6_out1_data;
	assign branch_6_in1_valid = phi_6_out1_valid;
	assign phi_6_out1_ready = branch_6_in1_ready;

	assign brCst_block4_clk = clk;
	assign brCst_block4_rst = rst;
	assign fork_12_in1_data = brCst_block4_out1_data;
	assign fork_12_in1_valid = brCst_block4_out1_valid;
	assign brCst_block4_out1_ready = fork_12_in1_ready;

	assign cst_3_clk = clk;
	assign cst_3_rst = rst;
	assign branch_5_in1_data = cst_3_out1_data;
	assign branch_5_in1_valid = cst_3_out1_valid;
	assign cst_3_out1_ready = branch_5_in1_ready;

	assign phi_n3_clk = clk;
	assign phi_n3_rst = rst;
	assign branch_7_in1_data = phi_n3_out1_data;
	assign branch_7_in1_valid = phi_n3_out1_valid;
	assign phi_n3_out1_ready = branch_7_in1_ready;

	assign branch_5_clk = clk;
	assign branch_5_rst = rst;
	assign phi_8_in2_data = branch_5_out1_data;
	assign phi_8_in2_valid = branch_5_out1_valid;
	assign branch_5_out1_ready = phi_8_in2_ready;
	assign sink_4_in1_data = branch_5_out2_data;
	assign sink_4_in1_valid = branch_5_out2_valid;
	assign branch_5_out2_ready = sink_4_in1_ready;

	assign branch_6_clk = clk;
	assign branch_6_rst = rst;
	assign phi_n6_in1_data = branch_6_out1_data;
	assign phi_n6_in1_valid = branch_6_out1_valid;
	assign branch_6_out1_ready = phi_n6_in1_ready;
	assign sink_5_in1_data = branch_6_out2_data;
	assign sink_5_in1_valid = branch_6_out2_valid;
	assign branch_6_out2_ready = sink_5_in1_ready;

	assign branch_7_clk = clk;
	assign branch_7_rst = rst;
	assign phi_n7_in1_data = branch_7_out1_data;
	assign phi_n7_in1_valid = branch_7_out1_valid;
	assign branch_7_out1_ready = phi_n7_in1_ready;
	assign sink_6_in1_data = branch_7_out2_data;
	assign sink_6_in1_valid = branch_7_out2_valid;
	assign branch_7_out2_ready = sink_6_in1_ready;

	assign fork_12_clk = clk;
	assign fork_12_rst = rst;
	assign branch_7_in2_data = fork_12_out1_data;
	assign branch_7_in2_valid = fork_12_out1_valid;
	assign fork_12_out1_ready = branch_7_in2_ready;
	assign branch_6_in2_data = fork_12_out2_data;
	assign branch_6_in2_valid = fork_12_out2_valid;
	assign fork_12_out2_ready = branch_6_in2_ready;
	assign branch_5_in2_data = fork_12_out3_data;
	assign branch_5_in2_valid = fork_12_out3_valid;
	assign fork_12_out3_ready = branch_5_in2_ready;
	assign branchC_17_in2_data = fork_12_out4_data;
	assign branchC_17_in2_valid = fork_12_out4_valid;
	assign fork_12_out4_ready = branchC_17_in2_ready;

	assign phiC_10_clk = clk;
	assign phiC_10_rst = rst;
	assign forkC_21_in1_data = phiC_10_out1_data;
	assign forkC_21_in1_valid = phiC_10_out1_valid;
	assign phiC_10_out1_ready = forkC_21_in1_ready;
	assign phi_6_in1_data = phiC_10_out2_data;
	assign phi_6_in1_valid = phiC_10_out2_valid;
	assign phiC_10_out2_ready = phi_6_in1_ready;

	assign forkC_21_clk = clk;
	assign forkC_21_rst = rst;
	assign cst_3_in1_data = forkC_21_out1_data;
	assign cst_3_in1_valid = forkC_21_out1_valid;
	assign forkC_21_out1_ready = cst_3_in1_ready;
	assign branchC_17_in1_data = forkC_21_out2_data;
	assign branchC_17_in1_valid = forkC_21_out2_valid;
	assign forkC_21_out2_ready = branchC_17_in1_ready;
	assign brCst_block4_in1_data = forkC_21_out3_data;
	assign brCst_block4_in1_valid = forkC_21_out3_valid;
	assign forkC_21_out3_ready = brCst_block4_in1_ready;

	assign branchC_17_clk = clk;
	assign branchC_17_rst = rst;
	assign phiC_11_in1_data = branchC_17_out1_data;
	assign phiC_11_in1_valid = branchC_17_out1_valid;
	assign branchC_17_out1_ready = phiC_11_in1_ready;
	assign sink_12_in1_data = branchC_17_out2_data;
	assign sink_12_in1_valid = branchC_17_out2_valid;
	assign branchC_17_out2_ready = sink_12_in1_ready;

	assign phi_8_clk = clk;
	assign phi_8_rst = rst;
	assign fork_2_in1_data = phi_8_out1_data;
	assign fork_2_in1_valid = phi_8_out1_valid;
	assign phi_8_out1_ready = fork_2_in1_ready;

	assign cst_4_clk = clk;
	assign cst_4_rst = rst;
	assign shl_9_in2_data = cst_4_out1_data;
	assign shl_9_in2_valid = cst_4_out1_valid;
	assign cst_4_out1_ready = shl_9_in2_ready;

	assign shl_9_clk = clk;
	assign shl_9_rst = rst;
	assign add_10_in1_data = shl_9_out1_data;
	assign add_10_in1_valid = shl_9_out1_valid;
	assign shl_9_out1_ready = add_10_in1_ready;

	assign add_10_clk = clk;
	assign add_10_rst = rst;
	assign load_13_in2_data = add_10_out1_data;
	assign load_13_in2_valid = add_10_out1_valid;
	assign add_10_out1_ready = load_13_in2_ready;

	assign load_13_clk = clk;
	assign load_13_rst = rst;
	assign sub_23_in1_data = load_13_out1_data;
	assign sub_23_in1_valid = load_13_out1_valid;
	assign load_13_out1_ready = sub_23_in1_ready;
	assign MC_A_in2_data = load_13_out2_data;
	assign MC_A_in2_valid = load_13_out2_valid;
	assign load_13_out2_ready = MC_A_in2_ready;

	assign load_16_clk = clk;
	assign load_16_rst = rst;
	assign mul_22_in1_data = load_16_out1_data;
	assign mul_22_in1_valid = load_16_out1_valid;
	assign load_16_out1_ready = mul_22_in1_ready;
	assign MC_c_in1_data = load_16_out2_data;
	assign MC_c_in1_valid = load_16_out2_valid;
	assign load_16_out2_ready = MC_c_in1_ready;

	assign cst_5_clk = clk;
	assign cst_5_rst = rst;
	assign shl_17_in2_data = cst_5_out1_data;
	assign shl_17_in2_valid = cst_5_out1_valid;
	assign cst_5_out1_ready = shl_17_in2_ready;

	assign shl_17_clk = clk;
	assign shl_17_rst = rst;
	assign add_18_in1_data = shl_17_out1_data;
	assign add_18_in1_valid = shl_17_out1_valid;
	assign shl_17_out1_ready = add_18_in1_ready;

	assign add_18_clk = clk;
	assign add_18_rst = rst;
	assign load_21_in2_data = add_18_out1_data;
	assign load_21_in2_valid = add_18_out1_valid;
	assign add_18_out1_ready = load_21_in2_ready;

	assign load_21_clk = clk;
	assign load_21_rst = rst;
	assign mul_22_in2_data = load_21_out1_data;
	assign mul_22_in2_valid = load_21_out1_valid;
	assign load_21_out1_ready = mul_22_in2_ready;
	assign MC_A_in3_data = load_21_out2_data;
	assign MC_A_in3_valid = load_21_out2_valid;
	assign load_21_out2_ready = MC_A_in3_ready;

	assign mul_22_clk = clk;
	assign mul_22_rst = rst;
	assign sub_23_in2_data = mul_22_out1_data;
	assign sub_23_in2_valid = mul_22_out1_valid;
	assign mul_22_out1_ready = sub_23_in2_ready;

	assign sub_23_clk = clk;
	assign sub_23_rst = rst;
	assign store_0_in1_data = sub_23_out1_data;
	assign store_0_in1_valid = sub_23_out1_valid;
	assign sub_23_out1_ready = store_0_in1_ready;

	assign cst_6_clk = clk;
	assign cst_6_rst = rst;
	assign shl_24_in2_data = cst_6_out1_data;
	assign shl_24_in2_valid = cst_6_out1_valid;
	assign cst_6_out1_ready = shl_24_in2_ready;

	assign shl_24_clk = clk;
	assign shl_24_rst = rst;
	assign add_25_in1_data = shl_24_out1_data;
	assign add_25_in1_valid = shl_24_out1_valid;
	assign shl_24_out1_ready = add_25_in1_ready;

	assign add_25_clk = clk;
	assign add_25_rst = rst;
	assign store_0_in2_data = add_25_out1_data;
	assign store_0_in2_valid = add_25_out1_valid;
	assign add_25_out1_ready = store_0_in2_ready;

	assign store_0_clk = clk;
	assign store_0_rst = rst;
	assign MC_A_in5_data = store_0_out1_data;
	assign MC_A_in5_valid = store_0_out1_valid;
	assign store_0_out1_ready = MC_A_in5_ready;
	assign MC_A_in4_data = store_0_out2_data;
	assign MC_A_in4_valid = store_0_out2_valid;
	assign store_0_out2_ready = MC_A_in4_ready;

	assign cst_7_clk = clk;
	assign cst_7_rst = rst;
	assign add_28_in2_data = cst_7_out1_data;
	assign add_28_in2_valid = cst_7_out1_valid;
	assign cst_7_out1_ready = add_28_in2_ready;

	assign add_28_clk = clk;
	assign add_28_rst = rst;
	assign fork_3_in1_data = add_28_out1_data;
	assign fork_3_in1_valid = add_28_out1_valid;
	assign add_28_out1_ready = fork_3_in1_ready;

	assign cst_8_clk = clk;
	assign cst_8_rst = rst;
	assign icmp_29_in2_data = cst_8_out1_data;
	assign icmp_29_in2_valid = cst_8_out1_valid;
	assign cst_8_out1_ready = icmp_29_in2_ready;

	assign icmp_29_clk = clk;
	assign icmp_29_rst = rst;
	assign fork_13_in1_data = icmp_29_out1_data;
	assign fork_13_in1_valid = icmp_29_out1_valid;
	assign icmp_29_out1_ready = fork_13_in1_ready;

	assign phi_n6_clk = clk;
	assign phi_n6_rst = rst;
	assign fork_7_in1_data = phi_n6_out1_data;
	assign fork_7_in1_valid = phi_n6_out1_valid;
	assign phi_n6_out1_ready = fork_7_in1_ready;

	assign phi_n7_clk = clk;
	assign phi_n7_rst = rst;
	assign fork_8_in1_data = phi_n7_out1_data;
	assign fork_8_in1_valid = phi_n7_out1_valid;
	assign phi_n7_out1_ready = fork_8_in1_ready;

	assign fork_2_clk = clk;
	assign fork_2_rst = rst;
	assign add_10_in2_data = fork_2_out1_data;
	assign add_10_in2_valid = fork_2_out1_valid;
	assign fork_2_out1_ready = add_10_in2_ready;
	assign add_18_in2_data = fork_2_out2_data;
	assign add_18_in2_valid = fork_2_out2_valid;
	assign fork_2_out2_ready = add_18_in2_ready;
	assign add_25_in2_data = fork_2_out3_data;
	assign add_25_in2_valid = fork_2_out3_valid;
	assign fork_2_out3_ready = add_25_in2_ready;
	assign add_28_in1_data = fork_2_out4_data;
	assign add_28_in1_valid = fork_2_out4_valid;
	assign fork_2_out4_ready = add_28_in1_ready;

	assign fork_3_clk = clk;
	assign fork_3_rst = rst;
	assign icmp_29_in1_data = fork_3_out1_data;
	assign icmp_29_in1_valid = fork_3_out1_valid;
	assign fork_3_out1_ready = icmp_29_in1_ready;
	assign branch_8_in1_data = fork_3_out2_data;
	assign branch_8_in1_valid = fork_3_out2_valid;
	assign fork_3_out2_ready = branch_8_in1_ready;

	assign fork_7_clk = clk;
	assign fork_7_rst = rst;
	assign shl_9_in1_data = fork_7_out1_data;
	assign shl_9_in1_valid = fork_7_out1_valid;
	assign fork_7_out1_ready = shl_9_in1_ready;
	assign shl_24_in1_data = fork_7_out2_data;
	assign shl_24_in1_valid = fork_7_out2_valid;
	assign fork_7_out2_ready = shl_24_in1_ready;
	assign branch_9_in1_data = fork_7_out3_data;
	assign branch_9_in1_valid = fork_7_out3_valid;
	assign fork_7_out3_ready = branch_9_in1_ready;

	assign fork_8_clk = clk;
	assign fork_8_rst = rst;
	assign load_16_in2_data = fork_8_out1_data;
	assign load_16_in2_valid = fork_8_out1_valid;
	assign fork_8_out1_ready = load_16_in2_ready;
	assign shl_17_in1_data = fork_8_out2_data;
	assign shl_17_in1_valid = fork_8_out2_valid;
	assign fork_8_out2_ready = shl_17_in1_ready;
	assign branch_10_in1_data = fork_8_out3_data;
	assign branch_10_in1_valid = fork_8_out3_valid;
	assign fork_8_out3_ready = branch_10_in1_ready;

	assign branch_8_clk = clk;
	assign branch_8_rst = rst;
	assign Buffer_100_in1_data = branch_8_out1_data;
	assign Buffer_100_in1_valid = branch_8_out1_valid;
	assign branch_8_out1_ready = Buffer_100_in1_ready;
	assign sink_7_in1_data = branch_8_out2_data;
	assign sink_7_in1_valid = branch_8_out2_valid;
	assign branch_8_out2_ready = sink_7_in1_ready;

	assign branch_9_clk = clk;
	assign branch_9_rst = rst;
	assign Buffer_101_in1_data = branch_9_out1_data;
	assign Buffer_101_in1_valid = branch_9_out1_valid;
	assign branch_9_out1_ready = Buffer_101_in1_ready;
	assign phi_n4_in1_data = branch_9_out2_data;
	assign phi_n4_in1_valid = branch_9_out2_valid;
	assign branch_9_out2_ready = phi_n4_in1_ready;

	assign branch_10_clk = clk;
	assign branch_10_rst = rst;
	assign Buffer_102_in1_data = branch_10_out1_data;
	assign Buffer_102_in1_valid = branch_10_out1_valid;
	assign branch_10_out1_ready = Buffer_102_in1_ready;
	assign phi_n5_in1_data = branch_10_out2_data;
	assign phi_n5_in1_valid = branch_10_out2_valid;
	assign branch_10_out2_ready = phi_n5_in1_ready;

	assign fork_13_clk = clk;
	assign fork_13_rst = rst;
	assign branch_10_in2_data = fork_13_out1_data;
	assign branch_10_in2_valid = fork_13_out1_valid;
	assign fork_13_out1_ready = branch_10_in2_ready;
	assign branch_9_in2_data = fork_13_out2_data;
	assign branch_9_in2_valid = fork_13_out2_valid;
	assign fork_13_out2_ready = branch_9_in2_ready;
	assign branch_8_in2_data = fork_13_out3_data;
	assign branch_8_in2_valid = fork_13_out3_valid;
	assign fork_13_out3_ready = branch_8_in2_ready;
	assign branchC_18_in2_data = fork_13_out4_data;
	assign branchC_18_in2_valid = fork_13_out4_valid;
	assign fork_13_out4_ready = branchC_18_in2_ready;

	assign cst_13_clk = clk;
	assign cst_13_rst = rst;
	assign MC_A_in1_data = cst_13_out1_data;
	assign MC_A_in1_valid = cst_13_out1_valid;
	assign cst_13_out1_ready = MC_A_in1_ready;

	assign phiC_11_clk = clk;
	assign phiC_11_rst = rst;
	assign forkC_22_in1_data = phiC_11_out1_data;
	assign forkC_22_in1_valid = phiC_11_out1_valid;
	assign phiC_11_out1_ready = forkC_22_in1_ready;
	assign phi_8_in1_data = phiC_11_out2_data;
	assign phi_8_in1_valid = phiC_11_out2_valid;
	assign phiC_11_out2_ready = phi_8_in1_ready;

	assign forkC_22_clk = clk;
	assign forkC_22_rst = rst;
	assign cst_13_in1_data = forkC_22_out1_data;
	assign cst_13_in1_valid = forkC_22_out1_valid;
	assign forkC_22_out1_ready = cst_13_in1_ready;
	assign branchC_18_in1_data = forkC_22_out2_data;
	assign branchC_18_in1_valid = forkC_22_out2_valid;
	assign forkC_22_out2_ready = branchC_18_in1_ready;

	assign branchC_18_clk = clk;
	assign branchC_18_rst = rst;
	assign Buffer_103_in1_data = branchC_18_out1_data;
	assign Buffer_103_in1_valid = branchC_18_out1_valid;
	assign branchC_18_out1_ready = Buffer_103_in1_ready;
	assign phiC_12_in1_data = branchC_18_out2_data;
	assign phiC_12_in1_valid = branchC_18_out2_valid;
	assign branchC_18_out2_ready = phiC_12_in1_ready;

	assign source_2_clk = clk;
	assign source_2_rst = rst;
	assign cst_4_in1_data = source_2_out1_data;
	assign cst_4_in1_valid = source_2_out1_valid;
	assign source_2_out1_ready = cst_4_in1_ready;

	assign source_3_clk = clk;
	assign source_3_rst = rst;
	assign cst_5_in1_data = source_3_out1_data;
	assign cst_5_in1_valid = source_3_out1_valid;
	assign source_3_out1_ready = cst_5_in1_ready;

	assign source_4_clk = clk;
	assign source_4_rst = rst;
	assign cst_6_in1_data = source_4_out1_data;
	assign cst_6_in1_valid = source_4_out1_valid;
	assign source_4_out1_ready = cst_6_in1_ready;

	assign source_5_clk = clk;
	assign source_5_rst = rst;
	assign cst_7_in1_data = source_5_out1_data;
	assign cst_7_in1_valid = source_5_out1_valid;
	assign source_5_out1_ready = cst_7_in1_ready;

	assign source_6_clk = clk;
	assign source_6_rst = rst;
	assign cst_8_in1_data = source_6_out1_data;
	assign cst_8_in1_valid = source_6_out1_valid;
	assign source_6_out1_ready = cst_8_in1_ready;

	assign phi_1_clk = clk;
	assign phi_1_rst = rst;
	assign fork_0_in1_data = phi_1_out1_data;
	assign fork_0_in1_valid = phi_1_out1_valid;
	assign phi_1_out1_ready = fork_0_in1_ready;

	assign cst_1_clk = clk;
	assign cst_1_rst = rst;
	assign add_2_in2_data = cst_1_out1_data;
	assign add_2_in2_valid = cst_1_out1_valid;
	assign cst_1_out1_ready = add_2_in2_ready;

	assign add_2_clk = clk;
	assign add_2_rst = rst;
	assign fork_1_in1_data = add_2_out1_data;
	assign fork_1_in1_valid = add_2_out1_valid;
	assign add_2_out1_ready = fork_1_in1_ready;

	assign cst_2_clk = clk;
	assign cst_2_rst = rst;
	assign icmp_3_in2_data = cst_2_out1_data;
	assign icmp_3_in2_valid = cst_2_out1_valid;
	assign cst_2_out1_ready = icmp_3_in2_ready;

	assign icmp_3_clk = clk;
	assign icmp_3_rst = rst;
	assign fork_10_in1_data = icmp_3_out1_data;
	assign fork_10_in1_valid = icmp_3_out1_valid;
	assign icmp_3_out1_ready = fork_10_in1_ready;

	assign fork_0_clk = clk;
	assign fork_0_rst = rst;
	assign add_2_in1_data = fork_0_out1_data;
	assign add_2_in1_valid = fork_0_out1_valid;
	assign fork_0_out1_ready = add_2_in1_ready;
	assign branch_1_in1_data = fork_0_out2_data;
	assign branch_1_in1_valid = fork_0_out2_valid;
	assign fork_0_out2_ready = branch_1_in1_ready;

	assign fork_1_clk = clk;
	assign fork_1_rst = rst;
	assign icmp_3_in1_data = fork_1_out1_data;
	assign icmp_3_in1_valid = fork_1_out1_valid;
	assign fork_1_out1_ready = icmp_3_in1_ready;
	assign branch_2_in1_data = fork_1_out2_data;
	assign branch_2_in1_valid = fork_1_out2_valid;
	assign fork_1_out2_ready = branch_2_in1_ready;

	assign branch_1_clk = clk;
	assign branch_1_rst = rst;
	assign phi_n2_in1_data = branch_1_out1_data;
	assign phi_n2_in1_valid = branch_1_out1_valid;
	assign branch_1_out1_ready = phi_n2_in1_ready;
	assign phi_n0_in1_data = branch_1_out2_data;
	assign phi_n0_in1_valid = branch_1_out2_valid;
	assign branch_1_out2_ready = phi_n0_in1_ready;

	assign branch_2_clk = clk;
	assign branch_2_rst = rst;
	assign phi_n1_in1_data = branch_2_out1_data;
	assign phi_n1_in1_valid = branch_2_out1_valid;
	assign branch_2_out1_ready = phi_n1_in1_ready;
	assign sink_1_in1_data = branch_2_out2_data;
	assign sink_1_in1_valid = branch_2_out2_valid;
	assign branch_2_out2_ready = sink_1_in1_ready;

	assign fork_10_clk = clk;
	assign fork_10_rst = rst;
	assign branch_2_in2_data = fork_10_out1_data;
	assign branch_2_in2_valid = fork_10_out1_valid;
	assign fork_10_out1_ready = branch_2_in2_ready;
	assign branch_1_in2_data = fork_10_out2_data;
	assign branch_1_in2_valid = fork_10_out2_valid;
	assign fork_10_out2_ready = branch_1_in2_ready;
	assign branchC_15_in2_data = fork_10_out3_data;
	assign branchC_15_in2_valid = fork_10_out3_valid;
	assign fork_10_out3_ready = branchC_15_in2_ready;

	assign phiC_8_clk = clk;
	assign phiC_8_rst = rst;
	assign branchC_15_in1_data = phiC_8_out1_data;
	assign branchC_15_in1_valid = phiC_8_out1_valid;
	assign phiC_8_out1_ready = branchC_15_in1_ready;
	assign phi_1_in1_data = phiC_8_out2_data;
	assign phi_1_in1_valid = phiC_8_out2_valid;
	assign phiC_8_out2_ready = phi_1_in1_ready;

	assign branchC_15_clk = clk;
	assign branchC_15_rst = rst;
	assign phiC_9_in1_data = branchC_15_out1_data;
	assign phiC_9_in1_valid = branchC_15_out1_valid;
	assign branchC_15_out1_ready = phiC_9_in1_ready;
	assign phiC_13_in1_data = branchC_15_out2_data;
	assign phiC_13_in1_valid = branchC_15_out2_valid;
	assign branchC_15_out2_ready = phiC_13_in1_ready;

	assign source_0_clk = clk;
	assign source_0_rst = rst;
	assign cst_1_in1_data = source_0_out1_data;
	assign cst_1_in1_valid = source_0_out1_valid;
	assign source_0_out1_ready = cst_1_in1_ready;

	assign source_1_clk = clk;
	assign source_1_rst = rst;
	assign cst_2_in1_data = source_1_out1_data;
	assign cst_2_in1_valid = source_1_out1_valid;
	assign source_1_out1_ready = cst_2_in1_ready;

	assign MC_A_clk = clk;
	assign MC_A_rst = rst;
	assign A_ce0 = A_we0;
	assign load_13_in1_data = MC_A_out1_data;
	assign load_13_in1_valid = MC_A_out1_valid;
	assign MC_A_out1_ready = load_13_in1_ready;
	assign load_21_in1_data = MC_A_out2_data;
	assign load_21_in1_valid = MC_A_out2_valid;
	assign MC_A_out2_ready = load_21_in1_ready;
	assign end_0_in1_data = MC_A_out3_data;
	assign end_0_in1_valid = MC_A_out3_valid;
	assign MC_A_out3_ready = end_0_in1_ready;

	assign MC_c_clk = clk;
	assign MC_c_rst = rst;
	assign c_ce0 = c_we0;
	assign MC_c_in2_valid = 0;
	assign MC_c_in2_data = 0;
	assign load_16_in1_data = MC_c_out1_data;
	assign load_16_in1_valid = MC_c_out1_valid;
	assign MC_c_out1_ready = load_16_in1_ready;
	assign end_0_in2_data = MC_c_out2_data;
	assign end_0_in2_valid = MC_c_out2_valid;
	assign MC_c_out2_ready = end_0_in2_ready;

	assign sink_0_clk = clk;
	assign sink_0_rst = rst;

	assign sink_1_clk = clk;
	assign sink_1_rst = rst;

	assign sink_2_clk = clk;
	assign sink_2_rst = rst;

	assign sink_3_clk = clk;
	assign sink_3_rst = rst;

	assign sink_4_clk = clk;
	assign sink_4_rst = rst;

	assign sink_5_clk = clk;
	assign sink_5_rst = rst;

	assign sink_6_clk = clk;
	assign sink_6_rst = rst;

	assign sink_7_clk = clk;
	assign sink_7_rst = rst;

	assign sink_8_clk = clk;
	assign sink_8_rst = rst;

	assign sink_9_clk = clk;
	assign sink_9_rst = rst;

	assign sink_10_clk = clk;
	assign sink_10_rst = rst;

	assign sink_11_clk = clk;
	assign sink_11_rst = rst;

	assign sink_12_clk = clk;
	assign sink_12_rst = rst;

	assign Buffer_100_clk = clk;
	assign Buffer_100_rst = rst;
	assign phi_8_in3_data = Buffer_100_out1_data;
	assign phi_8_in3_valid = Buffer_100_out1_valid;
	assign Buffer_100_out1_ready = phi_8_in3_ready;

	assign Buffer_101_clk = clk;
	assign Buffer_101_rst = rst;
	assign phi_n6_in2_data = Buffer_101_out1_data;
	assign phi_n6_in2_valid = Buffer_101_out1_valid;
	assign Buffer_101_out1_ready = phi_n6_in2_ready;

	assign Buffer_102_clk = clk;
	assign Buffer_102_rst = rst;
	assign phi_n7_in2_data = Buffer_102_out1_data;
	assign phi_n7_in2_valid = Buffer_102_out1_valid;
	assign Buffer_102_out1_ready = phi_n7_in2_ready;

	assign Buffer_103_clk = clk;
	assign Buffer_103_rst = rst;
	assign phiC_11_in2_data = Buffer_103_out1_data;
	assign phiC_11_in2_valid = Buffer_103_out1_valid;
	assign Buffer_103_out1_ready = phiC_11_in2_ready;

	assign Buffer_104_clk = clk;
	assign Buffer_104_rst = rst;
	assign phi_6_in3_data = Buffer_104_out1_data;
	assign phi_6_in3_valid = Buffer_104_out1_valid;
	assign Buffer_104_out1_ready = phi_6_in3_ready;

	assign Buffer_105_clk = clk;
	assign Buffer_105_rst = rst;
	assign phi_n3_in2_data = Buffer_105_out1_data;
	assign phi_n3_in2_valid = Buffer_105_out1_valid;
	assign Buffer_105_out1_ready = phi_n3_in2_ready;

	assign Buffer_106_clk = clk;
	assign Buffer_106_rst = rst;
	assign phiC_10_in2_data = Buffer_106_out1_data;
	assign phiC_10_in2_valid = Buffer_106_out1_valid;
	assign Buffer_106_out1_ready = phiC_10_in2_ready;

	assign Buffer_107_clk = clk;
	assign Buffer_107_rst = rst;
	assign phi_1_in3_data = Buffer_107_out1_data;
	assign phi_1_in3_valid = Buffer_107_out1_valid;
	assign Buffer_107_out1_ready = phi_1_in3_ready;

	assign Buffer_108_clk = clk;
	assign Buffer_108_rst = rst;
	assign phiC_8_in2_data = Buffer_108_out1_data;
	assign phiC_8_in2_valid = Buffer_108_out1_valid;
	assign Buffer_108_out1_ready = phiC_8_in2_ready;

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block1
		(.clk(brCst_block1_clk), .rst(brCst_block1_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block1_in1_valid}), .ready_in_bus({brCst_block1_in1_ready}), 
		.data_out_bus({brCst_block1_out1_data}), .valid_out_bus({brCst_block1_out1_valid}), .ready_out_bus({brCst_block1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_0
		(.clk(cst_0_clk), .rst(cst_0_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_0_in1_valid}), .ready_in_bus({cst_0_in1_ready}), 
		.data_out_bus({cst_0_out1_data}), .valid_out_bus({cst_0_out1_valid}), .ready_out_bus({cst_0_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_0
		(.clk(branch_0_clk), .rst(branch_0_rst),
		.data_in_bus({{branch_0_in2_data}, branch_0_in1_data}), .valid_in_bus({branch_0_in2_valid, branch_0_in1_valid}), .ready_in_bus({branch_0_in2_ready, branch_0_in1_ready}), 
		.data_out_bus({branch_0_out2_data, branch_0_out1_data}), .valid_out_bus({branch_0_out2_valid, branch_0_out1_valid}), .ready_out_bus({branch_0_out2_ready, branch_0_out1_ready}));

	start_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) start_node_start_0
		(.clk(start_0_clk), .rst(start_0_rst),
		.data_in_bus({start_0_in1_data}), .valid_in_bus({start_0_in1_valid}), .ready_in_bus({start_0_in1_ready}), 
		.data_out_bus({start_0_out1_data}), .valid_out_bus({start_0_out1_valid}), .ready_out_bus({start_0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_17
		(.clk(forkC_17_clk), .rst(forkC_17_rst),
		.data_in_bus({forkC_17_in1_data}), .valid_in_bus({forkC_17_in1_valid}), .ready_in_bus({forkC_17_in1_ready}), 
		.data_out_bus({forkC_17_out3_data, forkC_17_out2_data, forkC_17_out1_data}), .valid_out_bus({forkC_17_out3_valid, forkC_17_out2_valid, forkC_17_out1_valid}), .ready_out_bus({forkC_17_out3_ready, forkC_17_out2_ready, forkC_17_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_14
		(.clk(branchC_14_clk), .rst(branchC_14_rst),
		.data_in_bus({{branchC_14_in2_data}, branchC_14_in1_data}), .valid_in_bus({branchC_14_in2_valid, branchC_14_in1_valid}), .ready_in_bus({branchC_14_in2_ready, branchC_14_in1_ready}), 
		.data_out_bus({branchC_14_out2_data, branchC_14_out1_data}), .valid_out_bus({branchC_14_out2_valid, branchC_14_out1_valid}), .ready_out_bus({branchC_14_out2_ready, branchC_14_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_18
		(.clk(fork_18_clk), .rst(fork_18_rst),
		.data_in_bus({fork_18_in1_data}), .valid_in_bus({fork_18_in1_valid}), .ready_in_bus({fork_18_in1_ready}), 
		.data_out_bus({fork_18_out2_data, fork_18_out1_data}), .valid_out_bus({fork_18_out2_valid, fork_18_out1_valid}), .ready_out_bus({fork_18_out2_ready, fork_18_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block3
		(.clk(brCst_block3_clk), .rst(brCst_block3_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block3_in1_valid}), .ready_in_bus({brCst_block3_in1_ready}), 
		.data_out_bus({brCst_block3_out1_data}), .valid_out_bus({brCst_block3_out1_valid}), .ready_out_bus({brCst_block3_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n1
		(.clk(phi_n1_clk), .rst(phi_n1_rst),
		.data_in_bus({phi_n1_in1_data}), .valid_in_bus({phi_n1_in1_valid}), .ready_in_bus({phi_n1_in1_ready}), 
		.data_out_bus({phi_n1_out1_data}), .valid_out_bus({phi_n1_out1_valid}), .ready_out_bus({phi_n1_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n2
		(.clk(phi_n2_clk), .rst(phi_n2_rst),
		.data_in_bus({phi_n2_in1_data}), .valid_in_bus({phi_n2_in1_valid}), .ready_in_bus({phi_n2_in1_ready}), 
		.data_out_bus({phi_n2_out1_data}), .valid_out_bus({phi_n2_out1_valid}), .ready_out_bus({phi_n2_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_3
		(.clk(branch_3_clk), .rst(branch_3_rst),
		.data_in_bus({{5'b0, branch_3_in2_data}, branch_3_in1_data}), .valid_in_bus({branch_3_in2_valid, branch_3_in1_valid}), .ready_in_bus({branch_3_in2_ready, branch_3_in1_ready}), 
		.data_out_bus({branch_3_out2_data, branch_3_out1_data}), .valid_out_bus({branch_3_out2_valid, branch_3_out1_valid}), .ready_out_bus({branch_3_out2_ready, branch_3_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_4
		(.clk(branch_4_clk), .rst(branch_4_rst),
		.data_in_bus({{4'b0, branch_4_in2_data}, branch_4_in1_data}), .valid_in_bus({branch_4_in2_valid, branch_4_in1_valid}), .ready_in_bus({branch_4_in2_ready, branch_4_in1_ready}), 
		.data_out_bus({branch_4_out2_data, branch_4_out1_data}), .valid_out_bus({branch_4_out2_valid, branch_4_out1_valid}), .ready_out_bus({branch_4_out2_ready, branch_4_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_11
		(.clk(fork_11_clk), .rst(fork_11_rst),
		.data_in_bus({fork_11_in1_data}), .valid_in_bus({fork_11_in1_valid}), .ready_in_bus({fork_11_in1_ready}), 
		.data_out_bus({fork_11_out3_data, fork_11_out2_data, fork_11_out1_data}), .valid_out_bus({fork_11_out3_valid, fork_11_out2_valid, fork_11_out1_valid}), .ready_out_bus({fork_11_out3_ready, fork_11_out2_ready, fork_11_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_9
		(.clk(phiC_9_clk), .rst(phiC_9_rst),
		.data_in_bus({phiC_9_in1_data}), .valid_in_bus({phiC_9_in1_valid}), .ready_in_bus({phiC_9_in1_ready}), 
		.data_out_bus({phiC_9_out1_data}), .valid_out_bus({phiC_9_out1_valid}), .ready_out_bus({phiC_9_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_20
		(.clk(forkC_20_clk), .rst(forkC_20_rst),
		.data_in_bus({forkC_20_in1_data}), .valid_in_bus({forkC_20_in1_valid}), .ready_in_bus({forkC_20_in1_ready}), 
		.data_out_bus({forkC_20_out2_data, forkC_20_out1_data}), .valid_out_bus({forkC_20_out2_valid, forkC_20_out1_valid}), .ready_out_bus({forkC_20_out2_ready, forkC_20_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_16
		(.clk(branchC_16_clk), .rst(branchC_16_rst),
		.data_in_bus({{branchC_16_in2_data}, branchC_16_in1_data}), .valid_in_bus({branchC_16_in2_valid, branchC_16_in1_valid}), .ready_in_bus({branchC_16_in2_ready, branchC_16_in1_ready}), 
		.data_out_bus({branchC_16_out2_data, branchC_16_out1_data}), .valid_out_bus({branchC_16_out2_valid, branchC_16_out1_valid}), .ready_out_bus({branchC_16_out2_ready, branchC_16_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_9
		(.clk(cst_9_clk), .rst(cst_9_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_9_in1_valid}), .ready_in_bus({cst_9_in1_ready}), 
		.data_out_bus({cst_9_out1_data}), .valid_out_bus({cst_9_out1_valid}), .ready_out_bus({cst_9_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) add_op_add_31
		(.clk(add_31_clk), .rst(add_31_rst),
		.data_in_bus({add_31_in2_data, add_31_in1_data}), .valid_in_bus({add_31_in2_valid, add_31_in1_valid}), .ready_in_bus({add_31_in2_ready, add_31_in1_ready}), 
		.data_out_bus({add_31_out1_data}), .valid_out_bus({add_31_out1_valid}), .ready_out_bus({add_31_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) const_node_cst_10
		(.clk(cst_10_clk), .rst(cst_10_rst),
		.data_in_bus({4'd15}), .valid_in_bus({cst_10_in1_valid}), .ready_in_bus({cst_10_in1_ready}), 
		.data_out_bus({cst_10_out1_data}), .valid_out_bus({cst_10_out1_valid}), .ready_out_bus({cst_10_out1_ready}));

	icmp_slt_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_slt_op_icmp_32
		(.clk(icmp_32_clk), .rst(icmp_32_rst),
		.data_in_bus({icmp_32_in2_data, icmp_32_in1_data}), .valid_in_bus({icmp_32_in2_valid, icmp_32_in1_valid}), .ready_in_bus({icmp_32_in2_ready, icmp_32_in1_ready}), 
		.data_out_bus({icmp_32_out1_data}), .valid_out_bus({icmp_32_out1_valid}), .ready_out_bus({icmp_32_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n4
		(.clk(phi_n4_clk), .rst(phi_n4_rst),
		.data_in_bus({phi_n4_in1_data}), .valid_in_bus({phi_n4_in1_valid}), .ready_in_bus({phi_n4_in1_ready}), 
		.data_out_bus({phi_n4_out1_data}), .valid_out_bus({phi_n4_out1_valid}), .ready_out_bus({phi_n4_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n5
		(.clk(phi_n5_clk), .rst(phi_n5_rst),
		.data_in_bus({phi_n5_in1_data}), .valid_in_bus({phi_n5_in1_valid}), .ready_in_bus({phi_n5_in1_ready}), 
		.data_out_bus({phi_n5_out1_data}), .valid_out_bus({phi_n5_out1_valid}), .ready_out_bus({phi_n5_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_5
		(.clk(fork_5_clk), .rst(fork_5_rst),
		.data_in_bus({fork_5_in1_data}), .valid_in_bus({fork_5_in1_valid}), .ready_in_bus({fork_5_in1_ready}), 
		.data_out_bus({fork_5_out2_data, fork_5_out1_data}), .valid_out_bus({fork_5_out2_valid, fork_5_out1_valid}), .ready_out_bus({fork_5_out2_ready, fork_5_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_11
		(.clk(branch_11_clk), .rst(branch_11_rst),
		.data_in_bus({{4'b0, branch_11_in2_data}, branch_11_in1_data}), .valid_in_bus({branch_11_in2_valid, branch_11_in1_valid}), .ready_in_bus({branch_11_in2_ready, branch_11_in1_ready}), 
		.data_out_bus({branch_11_out2_data, branch_11_out1_data}), .valid_out_bus({branch_11_out2_valid, branch_11_out1_valid}), .ready_out_bus({branch_11_out2_ready, branch_11_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_12
		(.clk(branch_12_clk), .rst(branch_12_rst),
		.data_in_bus({{4'b0, branch_12_in2_data}, branch_12_in1_data}), .valid_in_bus({branch_12_in2_valid, branch_12_in1_valid}), .ready_in_bus({branch_12_in2_ready, branch_12_in1_ready}), 
		.data_out_bus({branch_12_out2_data, branch_12_out1_data}), .valid_out_bus({branch_12_out2_valid, branch_12_out1_valid}), .ready_out_bus({branch_12_out2_ready, branch_12_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_14
		(.clk(fork_14_clk), .rst(fork_14_rst),
		.data_in_bus({fork_14_in1_data}), .valid_in_bus({fork_14_in1_valid}), .ready_in_bus({fork_14_in1_ready}), 
		.data_out_bus({fork_14_out3_data, fork_14_out2_data, fork_14_out1_data}), .valid_out_bus({fork_14_out3_valid, fork_14_out2_valid, fork_14_out1_valid}), .ready_out_bus({fork_14_out3_ready, fork_14_out2_ready, fork_14_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_12
		(.clk(phiC_12_clk), .rst(phiC_12_rst),
		.data_in_bus({phiC_12_in1_data}), .valid_in_bus({phiC_12_in1_valid}), .ready_in_bus({phiC_12_in1_ready}), 
		.data_out_bus({phiC_12_out1_data}), .valid_out_bus({phiC_12_out1_valid}), .ready_out_bus({phiC_12_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_19
		(.clk(branchC_19_clk), .rst(branchC_19_rst),
		.data_in_bus({{branchC_19_in2_data}, branchC_19_in1_data}), .valid_in_bus({branchC_19_in2_valid, branchC_19_in1_valid}), .ready_in_bus({branchC_19_in2_ready, branchC_19_in1_ready}), 
		.data_out_bus({branchC_19_out2_data, branchC_19_out1_data}), .valid_out_bus({branchC_19_out2_valid, branchC_19_out1_valid}), .ready_out_bus({branchC_19_out2_ready, branchC_19_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_7
		(.clk(source_7_clk), .rst(source_7_rst),
		.data_out_bus({source_7_out1_data}), .valid_out_bus({source_7_out1_valid}), .ready_out_bus({source_7_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(4))source_node_source_8
		(.clk(source_8_clk), .rst(source_8_rst),
		.data_out_bus({source_8_out1_data}), .valid_out_bus({source_8_out1_valid}), .ready_out_bus({source_8_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_11
		(.clk(cst_11_clk), .rst(cst_11_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_11_in1_valid}), .ready_in_bus({cst_11_in1_ready}), 
		.data_out_bus({cst_11_out1_data}), .valid_out_bus({cst_11_out1_valid}), .ready_out_bus({cst_11_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) add_op_add_34
		(.clk(add_34_clk), .rst(add_34_rst),
		.data_in_bus({add_34_in2_data, add_34_in1_data}), .valid_in_bus({add_34_in2_valid, add_34_in1_valid}), .ready_in_bus({add_34_in2_ready, add_34_in1_ready}), 
		.data_out_bus({add_34_out1_data}), .valid_out_bus({add_34_out1_valid}), .ready_out_bus({add_34_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) const_node_cst_12
		(.clk(cst_12_clk), .rst(cst_12_rst),
		.data_in_bus({5'd16}), .valid_in_bus({cst_12_in1_valid}), .ready_in_bus({cst_12_in1_ready}), 
		.data_out_bus({cst_12_out1_data}), .valid_out_bus({cst_12_out1_valid}), .ready_out_bus({cst_12_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_35
		(.clk(icmp_35_clk), .rst(icmp_35_rst),
		.data_in_bus({icmp_35_in2_data, icmp_35_in1_data}), .valid_in_bus({icmp_35_in2_valid, icmp_35_in1_valid}), .ready_in_bus({icmp_35_in2_ready, icmp_35_in1_ready}), 
		.data_out_bus({icmp_35_out1_data}), .valid_out_bus({icmp_35_out1_valid}), .ready_out_bus({icmp_35_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n0
		(.clk(phi_n0_clk), .rst(phi_n0_rst),
		.data_in_bus({phi_n0_in2_data, phi_n0_in1_data}), .valid_in_bus({phi_n0_in2_valid, phi_n0_in1_valid}), .ready_in_bus({phi_n0_in2_ready, phi_n0_in1_ready}), 
		.data_out_bus({phi_n0_out1_data}), .valid_out_bus({phi_n0_out1_valid}), .ready_out_bus({phi_n0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_4
		(.clk(fork_4_clk), .rst(fork_4_rst),
		.data_in_bus({fork_4_in1_data}), .valid_in_bus({fork_4_in1_valid}), .ready_in_bus({fork_4_in1_ready}), 
		.data_out_bus({fork_4_out2_data, fork_4_out1_data}), .valid_out_bus({fork_4_out2_valid, fork_4_out1_valid}), .ready_out_bus({fork_4_out2_ready, fork_4_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_13
		(.clk(branch_13_clk), .rst(branch_13_rst),
		.data_in_bus({{4'b0, branch_13_in2_data}, branch_13_in1_data}), .valid_in_bus({branch_13_in2_valid, branch_13_in1_valid}), .ready_in_bus({branch_13_in2_ready, branch_13_in1_ready}), 
		.data_out_bus({branch_13_out2_data, branch_13_out1_data}), .valid_out_bus({branch_13_out2_valid, branch_13_out1_valid}), .ready_out_bus({branch_13_out2_ready, branch_13_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_13
		(.clk(phiC_13_clk), .rst(phiC_13_rst),
		.data_in_bus({phiC_13_in2_data, phiC_13_in1_data}), .valid_in_bus({phiC_13_in2_valid, phiC_13_in1_valid}), .ready_in_bus({phiC_13_in2_ready, phiC_13_in1_ready}), 
		.data_out_bus({phiC_13_out1_data}), .valid_out_bus({phiC_13_out1_valid}), .ready_out_bus({phiC_13_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_20
		(.clk(branchC_20_clk), .rst(branchC_20_rst),
		.data_in_bus({{branchC_20_in2_data}, branchC_20_in1_data}), .valid_in_bus({branchC_20_in2_valid, branchC_20_in1_valid}), .ready_in_bus({branchC_20_in2_ready, branchC_20_in1_ready}), 
		.data_out_bus({branchC_20_out2_data, branchC_20_out1_data}), .valid_out_bus({branchC_20_out2_valid, branchC_20_out1_valid}), .ready_out_bus({branchC_20_out2_ready, branchC_20_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_25
		(.clk(fork_25_clk), .rst(fork_25_rst),
		.data_in_bus({fork_25_in1_data}), .valid_in_bus({fork_25_in1_valid}), .ready_in_bus({fork_25_in1_ready}), 
		.data_out_bus({fork_25_out2_data, fork_25_out1_data}), .valid_out_bus({fork_25_out2_valid, fork_25_out1_valid}), .ready_out_bus({fork_25_out2_ready, fork_25_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_9
		(.clk(source_9_clk), .rst(source_9_rst),
		.data_out_bus({source_9_out1_data}), .valid_out_bus({source_9_out1_valid}), .ready_out_bus({source_9_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(5))source_node_source_10
		(.clk(source_10_clk), .rst(source_10_rst),
		.data_out_bus({source_10_out1_data}), .valid_out_bus({source_10_out1_valid}), .ready_out_bus({source_10_out1_ready}));

	ret_op #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) ret_op_ret_0
		(.clk(ret_0_clk), .rst(ret_0_rst),
		.data_in_bus({ret_0_in1_data}), .valid_in_bus({ret_0_in1_valid}), .ready_in_bus({ret_0_in1_ready}), 
		.data_out_bus({ret_0_out1_data}), .valid_out_bus({ret_0_out1_valid}), .ready_out_bus({ret_0_out1_ready}));

	end_node #(.INPUTS(1), .OUTPUTS(1), .MEMORY_INPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) end_node_end_0
		(.clk(end_0_clk), .rst(end_0_rst),
		.data_in_bus({end_0_in3_data}), .valid_in_bus({end_0_in3_valid}), .ready_in_bus({end_0_in3_ready}), .e_valid_bus({end_0_in2_valid, end_0_in1_valid}), .e_ready_bus({end_0_in2_ready, end_0_in1_ready}), 
		.data_out_bus({end_0_out1_data}), .valid_out_bus({end_0_out1_valid}), .ready_out_bus({end_0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_14
		(.clk(phiC_14_clk), .rst(phiC_14_rst),
		.data_in_bus({phiC_14_in1_data}), .valid_in_bus({phiC_14_in1_valid}), .ready_in_bus({phiC_14_in1_ready}), 
		.data_out_bus({phiC_14_out1_data}), .valid_out_bus({phiC_14_out1_valid}), .ready_out_bus({phiC_14_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5), .COND_SIZE(1)) mux_node_phi_6
		(.clk(phi_6_clk), .rst(phi_6_rst),
		.data_in_bus({{4'b0, phi_6_in1_data}, phi_6_in3_data, phi_6_in2_data}), .valid_in_bus({phi_6_in1_valid, phi_6_in3_valid, phi_6_in2_valid}), .ready_in_bus({phi_6_in1_ready, phi_6_in3_ready, phi_6_in2_ready}), 
		.data_out_bus({phi_6_out1_data}), .valid_out_bus({phi_6_out1_valid}), .ready_out_bus({phi_6_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block4
		(.clk(brCst_block4_clk), .rst(brCst_block4_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block4_in1_valid}), .ready_in_bus({brCst_block4_in1_ready}), 
		.data_out_bus({brCst_block4_out1_data}), .valid_out_bus({brCst_block4_out1_valid}), .ready_out_bus({brCst_block4_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_3
		(.clk(cst_3_clk), .rst(cst_3_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_3_in1_valid}), .ready_in_bus({cst_3_in1_ready}), 
		.data_out_bus({cst_3_out1_data}), .valid_out_bus({cst_3_out1_valid}), .ready_out_bus({cst_3_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n3
		(.clk(phi_n3_clk), .rst(phi_n3_rst),
		.data_in_bus({phi_n3_in2_data, phi_n3_in1_data}), .valid_in_bus({phi_n3_in2_valid, phi_n3_in1_valid}), .ready_in_bus({phi_n3_in2_ready, phi_n3_in1_ready}), 
		.data_out_bus({phi_n3_out1_data}), .valid_out_bus({phi_n3_out1_valid}), .ready_out_bus({phi_n3_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_5
		(.clk(branch_5_clk), .rst(branch_5_rst),
		.data_in_bus({{branch_5_in2_data}, branch_5_in1_data}), .valid_in_bus({branch_5_in2_valid, branch_5_in1_valid}), .ready_in_bus({branch_5_in2_ready, branch_5_in1_ready}), 
		.data_out_bus({branch_5_out2_data, branch_5_out1_data}), .valid_out_bus({branch_5_out2_valid, branch_5_out1_valid}), .ready_out_bus({branch_5_out2_ready, branch_5_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_6
		(.clk(branch_6_clk), .rst(branch_6_rst),
		.data_in_bus({{4'b0, branch_6_in2_data}, branch_6_in1_data}), .valid_in_bus({branch_6_in2_valid, branch_6_in1_valid}), .ready_in_bus({branch_6_in2_ready, branch_6_in1_ready}), 
		.data_out_bus({branch_6_out2_data, branch_6_out1_data}), .valid_out_bus({branch_6_out2_valid, branch_6_out1_valid}), .ready_out_bus({branch_6_out2_ready, branch_6_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_7
		(.clk(branch_7_clk), .rst(branch_7_rst),
		.data_in_bus({{4'b0, branch_7_in2_data}, branch_7_in1_data}), .valid_in_bus({branch_7_in2_valid, branch_7_in1_valid}), .ready_in_bus({branch_7_in2_ready, branch_7_in1_ready}), 
		.data_out_bus({branch_7_out2_data, branch_7_out1_data}), .valid_out_bus({branch_7_out2_valid, branch_7_out1_valid}), .ready_out_bus({branch_7_out2_ready, branch_7_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_12
		(.clk(fork_12_clk), .rst(fork_12_rst),
		.data_in_bus({fork_12_in1_data}), .valid_in_bus({fork_12_in1_valid}), .ready_in_bus({fork_12_in1_ready}), 
		.data_out_bus({fork_12_out4_data, fork_12_out3_data, fork_12_out2_data, fork_12_out1_data}), .valid_out_bus({fork_12_out4_valid, fork_12_out3_valid, fork_12_out2_valid, fork_12_out1_valid}), .ready_out_bus({fork_12_out4_ready, fork_12_out3_ready, fork_12_out2_ready, fork_12_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_10
		(.clk(phiC_10_clk), .rst(phiC_10_rst),
		.data_in_bus({phiC_10_in2_data, phiC_10_in1_data}), .valid_in_bus({phiC_10_in2_valid, phiC_10_in1_valid}), .ready_in_bus({phiC_10_in2_ready, phiC_10_in1_ready}), 
		.data_out_bus({phiC_10_out2_data, phiC_10_out1_data}), .valid_out_bus({phiC_10_out2_valid, phiC_10_out1_valid}), .ready_out_bus({phiC_10_out2_ready, phiC_10_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_21
		(.clk(forkC_21_clk), .rst(forkC_21_rst),
		.data_in_bus({forkC_21_in1_data}), .valid_in_bus({forkC_21_in1_valid}), .ready_in_bus({forkC_21_in1_ready}), 
		.data_out_bus({forkC_21_out3_data, forkC_21_out2_data, forkC_21_out1_data}), .valid_out_bus({forkC_21_out3_valid, forkC_21_out2_valid, forkC_21_out1_valid}), .ready_out_bus({forkC_21_out3_ready, forkC_21_out2_ready, forkC_21_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_17
		(.clk(branchC_17_clk), .rst(branchC_17_rst),
		.data_in_bus({{branchC_17_in2_data}, branchC_17_in1_data}), .valid_in_bus({branchC_17_in2_valid, branchC_17_in1_valid}), .ready_in_bus({branchC_17_in2_ready, branchC_17_in1_ready}), 
		.data_out_bus({branchC_17_out2_data, branchC_17_out1_data}), .valid_out_bus({branchC_17_out2_valid, branchC_17_out1_valid}), .ready_out_bus({branchC_17_out2_ready, branchC_17_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5), .COND_SIZE(1)) mux_node_phi_8
		(.clk(phi_8_clk), .rst(phi_8_rst),
		.data_in_bus({{4'b0, phi_8_in1_data}, phi_8_in3_data, phi_8_in2_data}), .valid_in_bus({phi_8_in1_valid, phi_8_in3_valid, phi_8_in2_valid}), .ready_in_bus({phi_8_in1_ready, phi_8_in3_ready, phi_8_in2_ready}), 
		.data_out_bus({phi_8_out1_data}), .valid_out_bus({phi_8_out1_valid}), .ready_out_bus({phi_8_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_4
		(.clk(cst_4_clk), .rst(cst_4_rst),
		.data_in_bus({3'd4}), .valid_in_bus({cst_4_in1_valid}), .ready_in_bus({cst_4_in1_ready}), 
		.data_out_bus({cst_4_out1_data}), .valid_out_bus({cst_4_out1_valid}), .ready_out_bus({cst_4_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(9), .DATA_OUT_SIZE(9)) shl_op_shl_9
		(.clk(shl_9_clk), .rst(shl_9_rst),
		.data_in_bus({shl_9_in2_data, shl_9_in1_data}), .valid_in_bus({shl_9_in2_valid, shl_9_in1_valid}), .ready_in_bus({shl_9_in2_ready, shl_9_in1_ready}), 
		.data_out_bus({shl_9_out1_data}), .valid_out_bus({shl_9_out1_valid}), .ready_out_bus({shl_9_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) add_op_add_10
		(.clk(add_10_clk), .rst(add_10_rst),
		.data_in_bus({add_10_in2_data, add_10_in1_data}), .valid_in_bus({add_10_in2_valid, add_10_in1_valid}), .ready_in_bus({add_10_in2_ready, add_10_in1_ready}), 
		.data_out_bus({add_10_out1_data}), .valid_out_bus({add_10_out1_valid}), .ready_out_bus({add_10_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(10), .DATA_SIZE(32)) mc_load_op_load_13
		(.clk(load_13_clk), .rst(load_13_rst),
		.data_in_bus({load_13_in1_data}), .address_in_bus({load_13_in2_data}), .valid_in_bus({load_13_in2_valid, load_13_in1_valid}), .ready_in_bus({load_13_in2_ready, load_13_in1_ready}), 
		.data_out_bus({load_13_out1_data}), .address_out_bus({load_13_out2_data}), .valid_out_bus({load_13_out2_valid, load_13_out1_valid}), .ready_out_bus({load_13_out2_ready, load_13_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(5), .DATA_SIZE(32)) mc_load_op_load_16
		(.clk(load_16_clk), .rst(load_16_rst),
		.data_in_bus({load_16_in1_data}), .address_in_bus({load_16_in2_data}), .valid_in_bus({load_16_in2_valid, load_16_in1_valid}), .ready_in_bus({load_16_in2_ready, load_16_in1_ready}), 
		.data_out_bus({load_16_out1_data}), .address_out_bus({load_16_out2_data}), .valid_out_bus({load_16_out2_valid, load_16_out1_valid}), .ready_out_bus({load_16_out2_ready, load_16_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_5
		(.clk(cst_5_clk), .rst(cst_5_rst),
		.data_in_bus({3'd4}), .valid_in_bus({cst_5_in1_valid}), .ready_in_bus({cst_5_in1_ready}), 
		.data_out_bus({cst_5_out1_data}), .valid_out_bus({cst_5_out1_valid}), .ready_out_bus({cst_5_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(9), .DATA_OUT_SIZE(9)) shl_op_shl_17
		(.clk(shl_17_clk), .rst(shl_17_rst),
		.data_in_bus({shl_17_in2_data, shl_17_in1_data}), .valid_in_bus({shl_17_in2_valid, shl_17_in1_valid}), .ready_in_bus({shl_17_in2_ready, shl_17_in1_ready}), 
		.data_out_bus({shl_17_out1_data}), .valid_out_bus({shl_17_out1_valid}), .ready_out_bus({shl_17_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) add_op_add_18
		(.clk(add_18_clk), .rst(add_18_rst),
		.data_in_bus({add_18_in2_data, add_18_in1_data}), .valid_in_bus({add_18_in2_valid, add_18_in1_valid}), .ready_in_bus({add_18_in2_ready, add_18_in1_ready}), 
		.data_out_bus({add_18_out1_data}), .valid_out_bus({add_18_out1_valid}), .ready_out_bus({add_18_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(10), .DATA_SIZE(32)) mc_load_op_load_21
		(.clk(load_21_clk), .rst(load_21_rst),
		.data_in_bus({load_21_in1_data}), .address_in_bus({load_21_in2_data}), .valid_in_bus({load_21_in2_valid, load_21_in1_valid}), .ready_in_bus({load_21_in2_ready, load_21_in1_ready}), 
		.data_out_bus({load_21_out1_data}), .address_out_bus({load_21_out2_data}), .valid_out_bus({load_21_out2_valid, load_21_out1_valid}), .ready_out_bus({load_21_out2_ready, load_21_out1_ready}));

	mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(16), .DATA_OUT_SIZE(32)) mul_op_mul_22
		(.clk(mul_22_clk), .rst(mul_22_rst),
		.data_in_bus({mul_22_in2_data, mul_22_in1_data}), .valid_in_bus({mul_22_in2_valid, mul_22_in1_valid}), .ready_in_bus({mul_22_in2_ready, mul_22_in1_ready}), 
		.data_out_bus({mul_22_out1_data}), .valid_out_bus({mul_22_out1_valid}), .ready_out_bus({mul_22_out1_ready}));

	sub_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) sub_op_sub_23
		(.clk(sub_23_clk), .rst(sub_23_rst),
		.data_in_bus({sub_23_in2_data, sub_23_in1_data}), .valid_in_bus({sub_23_in2_valid, sub_23_in1_valid}), .ready_in_bus({sub_23_in2_ready, sub_23_in1_ready}), 
		.data_out_bus({sub_23_out1_data}), .valid_out_bus({sub_23_out1_valid}), .ready_out_bus({sub_23_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_6
		(.clk(cst_6_clk), .rst(cst_6_rst),
		.data_in_bus({3'd4}), .valid_in_bus({cst_6_in1_valid}), .ready_in_bus({cst_6_in1_ready}), 
		.data_out_bus({cst_6_out1_data}), .valid_out_bus({cst_6_out1_valid}), .ready_out_bus({cst_6_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(9), .DATA_OUT_SIZE(9)) shl_op_shl_24
		(.clk(shl_24_clk), .rst(shl_24_rst),
		.data_in_bus({shl_24_in2_data, shl_24_in1_data}), .valid_in_bus({shl_24_in2_valid, shl_24_in1_valid}), .ready_in_bus({shl_24_in2_ready, shl_24_in1_ready}), 
		.data_out_bus({shl_24_out1_data}), .valid_out_bus({shl_24_out1_valid}), .ready_out_bus({shl_24_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) add_op_add_25
		(.clk(add_25_clk), .rst(add_25_rst),
		.data_in_bus({add_25_in2_data, add_25_in1_data}), .valid_in_bus({add_25_in2_valid, add_25_in1_valid}), .ready_in_bus({add_25_in2_ready, add_25_in1_ready}), 
		.data_out_bus({add_25_out1_data}), .valid_out_bus({add_25_out1_valid}), .ready_out_bus({add_25_out1_ready}));

	mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(10), .DATA_SIZE(32)) mc_store_op_store_0
		(.clk(store_0_clk), .rst(store_0_rst),
		.data_in_bus({store_0_in1_data}), .address_in_bus({store_0_in2_data}), .valid_in_bus({store_0_in2_valid, store_0_in1_valid}), .ready_in_bus({store_0_in2_ready, store_0_in1_ready}), 
		.data_out_bus({store_0_out1_data}), .address_out_bus({store_0_out2_data}), .valid_out_bus({store_0_out2_valid, store_0_out1_valid}), .ready_out_bus({store_0_out2_ready, store_0_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_7
		(.clk(cst_7_clk), .rst(cst_7_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_7_in1_valid}), .ready_in_bus({cst_7_in1_ready}), 
		.data_out_bus({cst_7_out1_data}), .valid_out_bus({cst_7_out1_valid}), .ready_out_bus({cst_7_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) add_op_add_28
		(.clk(add_28_clk), .rst(add_28_rst),
		.data_in_bus({add_28_in2_data, add_28_in1_data}), .valid_in_bus({add_28_in2_valid, add_28_in1_valid}), .ready_in_bus({add_28_in2_ready, add_28_in1_ready}), 
		.data_out_bus({add_28_out1_data}), .valid_out_bus({add_28_out1_valid}), .ready_out_bus({add_28_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) const_node_cst_8
		(.clk(cst_8_clk), .rst(cst_8_rst),
		.data_in_bus({5'd16}), .valid_in_bus({cst_8_in1_valid}), .ready_in_bus({cst_8_in1_ready}), 
		.data_out_bus({cst_8_out1_data}), .valid_out_bus({cst_8_out1_valid}), .ready_out_bus({cst_8_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_29
		(.clk(icmp_29_clk), .rst(icmp_29_rst),
		.data_in_bus({icmp_29_in2_data, icmp_29_in1_data}), .valid_in_bus({icmp_29_in2_valid, icmp_29_in1_valid}), .ready_in_bus({icmp_29_in2_ready, icmp_29_in1_ready}), 
		.data_out_bus({icmp_29_out1_data}), .valid_out_bus({icmp_29_out1_valid}), .ready_out_bus({icmp_29_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n6
		(.clk(phi_n6_clk), .rst(phi_n6_rst),
		.data_in_bus({phi_n6_in2_data, phi_n6_in1_data}), .valid_in_bus({phi_n6_in2_valid, phi_n6_in1_valid}), .ready_in_bus({phi_n6_in2_ready, phi_n6_in1_ready}), 
		.data_out_bus({phi_n6_out1_data}), .valid_out_bus({phi_n6_out1_valid}), .ready_out_bus({phi_n6_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n7
		(.clk(phi_n7_clk), .rst(phi_n7_rst),
		.data_in_bus({phi_n7_in2_data, phi_n7_in1_data}), .valid_in_bus({phi_n7_in2_valid, phi_n7_in1_valid}), .ready_in_bus({phi_n7_in2_ready, phi_n7_in1_ready}), 
		.data_out_bus({phi_n7_out1_data}), .valid_out_bus({phi_n7_out1_valid}), .ready_out_bus({phi_n7_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_2
		(.clk(fork_2_clk), .rst(fork_2_rst),
		.data_in_bus({fork_2_in1_data}), .valid_in_bus({fork_2_in1_valid}), .ready_in_bus({fork_2_in1_ready}), 
		.data_out_bus({fork_2_out4_data, fork_2_out3_data, fork_2_out2_data, fork_2_out1_data}), .valid_out_bus({fork_2_out4_valid, fork_2_out3_valid, fork_2_out2_valid, fork_2_out1_valid}), .ready_out_bus({fork_2_out4_ready, fork_2_out3_ready, fork_2_out2_ready, fork_2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_3
		(.clk(fork_3_clk), .rst(fork_3_rst),
		.data_in_bus({fork_3_in1_data}), .valid_in_bus({fork_3_in1_valid}), .ready_in_bus({fork_3_in1_ready}), 
		.data_out_bus({fork_3_out2_data, fork_3_out1_data}), .valid_out_bus({fork_3_out2_valid, fork_3_out1_valid}), .ready_out_bus({fork_3_out2_ready, fork_3_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_7
		(.clk(fork_7_clk), .rst(fork_7_rst),
		.data_in_bus({fork_7_in1_data}), .valid_in_bus({fork_7_in1_valid}), .ready_in_bus({fork_7_in1_ready}), 
		.data_out_bus({fork_7_out3_data, fork_7_out2_data, fork_7_out1_data}), .valid_out_bus({fork_7_out3_valid, fork_7_out2_valid, fork_7_out1_valid}), .ready_out_bus({fork_7_out3_ready, fork_7_out2_ready, fork_7_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_8
		(.clk(fork_8_clk), .rst(fork_8_rst),
		.data_in_bus({fork_8_in1_data}), .valid_in_bus({fork_8_in1_valid}), .ready_in_bus({fork_8_in1_ready}), 
		.data_out_bus({fork_8_out3_data, fork_8_out2_data, fork_8_out1_data}), .valid_out_bus({fork_8_out3_valid, fork_8_out2_valid, fork_8_out1_valid}), .ready_out_bus({fork_8_out3_ready, fork_8_out2_ready, fork_8_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_8
		(.clk(branch_8_clk), .rst(branch_8_rst),
		.data_in_bus({{4'b0, branch_8_in2_data}, branch_8_in1_data}), .valid_in_bus({branch_8_in2_valid, branch_8_in1_valid}), .ready_in_bus({branch_8_in2_ready, branch_8_in1_ready}), 
		.data_out_bus({branch_8_out2_data, branch_8_out1_data}), .valid_out_bus({branch_8_out2_valid, branch_8_out1_valid}), .ready_out_bus({branch_8_out2_ready, branch_8_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_9
		(.clk(branch_9_clk), .rst(branch_9_rst),
		.data_in_bus({{4'b0, branch_9_in2_data}, branch_9_in1_data}), .valid_in_bus({branch_9_in2_valid, branch_9_in1_valid}), .ready_in_bus({branch_9_in2_ready, branch_9_in1_ready}), 
		.data_out_bus({branch_9_out2_data, branch_9_out1_data}), .valid_out_bus({branch_9_out2_valid, branch_9_out1_valid}), .ready_out_bus({branch_9_out2_ready, branch_9_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_10
		(.clk(branch_10_clk), .rst(branch_10_rst),
		.data_in_bus({{4'b0, branch_10_in2_data}, branch_10_in1_data}), .valid_in_bus({branch_10_in2_valid, branch_10_in1_valid}), .ready_in_bus({branch_10_in2_ready, branch_10_in1_ready}), 
		.data_out_bus({branch_10_out2_data, branch_10_out1_data}), .valid_out_bus({branch_10_out2_valid, branch_10_out1_valid}), .ready_out_bus({branch_10_out2_ready, branch_10_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_13
		(.clk(fork_13_clk), .rst(fork_13_rst),
		.data_in_bus({fork_13_in1_data}), .valid_in_bus({fork_13_in1_valid}), .ready_in_bus({fork_13_in1_ready}), 
		.data_out_bus({fork_13_out4_data, fork_13_out3_data, fork_13_out2_data, fork_13_out1_data}), .valid_out_bus({fork_13_out4_valid, fork_13_out3_valid, fork_13_out2_valid, fork_13_out1_valid}), .ready_out_bus({fork_13_out4_ready, fork_13_out3_ready, fork_13_out2_ready, fork_13_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_13
		(.clk(cst_13_clk), .rst(cst_13_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_13_in1_valid}), .ready_in_bus({cst_13_in1_ready}), 
		.data_out_bus({cst_13_out1_data}), .valid_out_bus({cst_13_out1_valid}), .ready_out_bus({cst_13_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_11
		(.clk(phiC_11_clk), .rst(phiC_11_rst),
		.data_in_bus({phiC_11_in2_data, phiC_11_in1_data}), .valid_in_bus({phiC_11_in2_valid, phiC_11_in1_valid}), .ready_in_bus({phiC_11_in2_ready, phiC_11_in1_ready}), 
		.data_out_bus({phiC_11_out2_data, phiC_11_out1_data}), .valid_out_bus({phiC_11_out2_valid, phiC_11_out1_valid}), .ready_out_bus({phiC_11_out2_ready, phiC_11_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_22
		(.clk(forkC_22_clk), .rst(forkC_22_rst),
		.data_in_bus({forkC_22_in1_data}), .valid_in_bus({forkC_22_in1_valid}), .ready_in_bus({forkC_22_in1_ready}), 
		.data_out_bus({forkC_22_out2_data, forkC_22_out1_data}), .valid_out_bus({forkC_22_out2_valid, forkC_22_out1_valid}), .ready_out_bus({forkC_22_out2_ready, forkC_22_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_18
		(.clk(branchC_18_clk), .rst(branchC_18_rst),
		.data_in_bus({{branchC_18_in2_data}, branchC_18_in1_data}), .valid_in_bus({branchC_18_in2_valid, branchC_18_in1_valid}), .ready_in_bus({branchC_18_in2_ready, branchC_18_in1_ready}), 
		.data_out_bus({branchC_18_out2_data, branchC_18_out1_data}), .valid_out_bus({branchC_18_out2_valid, branchC_18_out1_valid}), .ready_out_bus({branchC_18_out2_ready, branchC_18_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_2
		(.clk(source_2_clk), .rst(source_2_rst),
		.data_out_bus({source_2_out1_data}), .valid_out_bus({source_2_out1_valid}), .ready_out_bus({source_2_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_3
		(.clk(source_3_clk), .rst(source_3_rst),
		.data_out_bus({source_3_out1_data}), .valid_out_bus({source_3_out1_valid}), .ready_out_bus({source_3_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_4
		(.clk(source_4_clk), .rst(source_4_rst),
		.data_out_bus({source_4_out1_data}), .valid_out_bus({source_4_out1_valid}), .ready_out_bus({source_4_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_5
		(.clk(source_5_clk), .rst(source_5_rst),
		.data_out_bus({source_5_out1_data}), .valid_out_bus({source_5_out1_valid}), .ready_out_bus({source_5_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(5))source_node_source_6
		(.clk(source_6_clk), .rst(source_6_rst),
		.data_out_bus({source_6_out1_data}), .valid_out_bus({source_6_out1_valid}), .ready_out_bus({source_6_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5), .COND_SIZE(1)) mux_node_phi_1
		(.clk(phi_1_clk), .rst(phi_1_rst),
		.data_in_bus({{4'b0, phi_1_in1_data}, phi_1_in3_data, phi_1_in2_data}), .valid_in_bus({phi_1_in1_valid, phi_1_in3_valid, phi_1_in2_valid}), .ready_in_bus({phi_1_in1_ready, phi_1_in3_ready, phi_1_in2_ready}), 
		.data_out_bus({phi_1_out1_data}), .valid_out_bus({phi_1_out1_valid}), .ready_out_bus({phi_1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_1
		(.clk(cst_1_clk), .rst(cst_1_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_1_in1_valid}), .ready_in_bus({cst_1_in1_ready}), 
		.data_out_bus({cst_1_out1_data}), .valid_out_bus({cst_1_out1_valid}), .ready_out_bus({cst_1_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_2
		(.clk(add_2_clk), .rst(add_2_rst),
		.data_in_bus({add_2_in2_data, add_2_in1_data}), .valid_in_bus({add_2_in2_valid, add_2_in1_valid}), .ready_in_bus({add_2_in2_ready, add_2_in1_ready}), 
		.data_out_bus({add_2_out1_data}), .valid_out_bus({add_2_out1_valid}), .ready_out_bus({add_2_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) const_node_cst_2
		(.clk(cst_2_clk), .rst(cst_2_rst),
		.data_in_bus({5'd16}), .valid_in_bus({cst_2_in1_valid}), .ready_in_bus({cst_2_in1_ready}), 
		.data_out_bus({cst_2_out1_data}), .valid_out_bus({cst_2_out1_valid}), .ready_out_bus({cst_2_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_3
		(.clk(icmp_3_clk), .rst(icmp_3_rst),
		.data_in_bus({icmp_3_in2_data, icmp_3_in1_data}), .valid_in_bus({icmp_3_in2_valid, icmp_3_in1_valid}), .ready_in_bus({icmp_3_in2_ready, icmp_3_in1_ready}), 
		.data_out_bus({icmp_3_out1_data}), .valid_out_bus({icmp_3_out1_valid}), .ready_out_bus({icmp_3_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_0
		(.clk(fork_0_clk), .rst(fork_0_rst),
		.data_in_bus({fork_0_in1_data}), .valid_in_bus({fork_0_in1_valid}), .ready_in_bus({fork_0_in1_ready}), 
		.data_out_bus({fork_0_out2_data, fork_0_out1_data}), .valid_out_bus({fork_0_out2_valid, fork_0_out1_valid}), .ready_out_bus({fork_0_out2_ready, fork_0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_1
		(.clk(fork_1_clk), .rst(fork_1_rst),
		.data_in_bus({fork_1_in1_data}), .valid_in_bus({fork_1_in1_valid}), .ready_in_bus({fork_1_in1_ready}), 
		.data_out_bus({fork_1_out2_data, fork_1_out1_data}), .valid_out_bus({fork_1_out2_valid, fork_1_out1_valid}), .ready_out_bus({fork_1_out2_ready, fork_1_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_1
		(.clk(branch_1_clk), .rst(branch_1_rst),
		.data_in_bus({{4'b0, branch_1_in2_data}, branch_1_in1_data}), .valid_in_bus({branch_1_in2_valid, branch_1_in1_valid}), .ready_in_bus({branch_1_in2_ready, branch_1_in1_ready}), 
		.data_out_bus({branch_1_out2_data, branch_1_out1_data}), .valid_out_bus({branch_1_out2_valid, branch_1_out1_valid}), .ready_out_bus({branch_1_out2_ready, branch_1_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_2
		(.clk(branch_2_clk), .rst(branch_2_rst),
		.data_in_bus({{5'b0, branch_2_in2_data}, branch_2_in1_data}), .valid_in_bus({branch_2_in2_valid, branch_2_in1_valid}), .ready_in_bus({branch_2_in2_ready, branch_2_in1_ready}), 
		.data_out_bus({branch_2_out2_data, branch_2_out1_data}), .valid_out_bus({branch_2_out2_valid, branch_2_out1_valid}), .ready_out_bus({branch_2_out2_ready, branch_2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_10
		(.clk(fork_10_clk), .rst(fork_10_rst),
		.data_in_bus({fork_10_in1_data}), .valid_in_bus({fork_10_in1_valid}), .ready_in_bus({fork_10_in1_ready}), 
		.data_out_bus({fork_10_out3_data, fork_10_out2_data, fork_10_out1_data}), .valid_out_bus({fork_10_out3_valid, fork_10_out2_valid, fork_10_out1_valid}), .ready_out_bus({fork_10_out3_ready, fork_10_out2_ready, fork_10_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_8
		(.clk(phiC_8_clk), .rst(phiC_8_rst),
		.data_in_bus({phiC_8_in2_data, phiC_8_in1_data}), .valid_in_bus({phiC_8_in2_valid, phiC_8_in1_valid}), .ready_in_bus({phiC_8_in2_ready, phiC_8_in1_ready}), 
		.data_out_bus({phiC_8_out2_data, phiC_8_out1_data}), .valid_out_bus({phiC_8_out2_valid, phiC_8_out1_valid}), .ready_out_bus({phiC_8_out2_ready, phiC_8_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_15
		(.clk(branchC_15_clk), .rst(branchC_15_rst),
		.data_in_bus({{branchC_15_in2_data}, branchC_15_in1_data}), .valid_in_bus({branchC_15_in2_valid, branchC_15_in1_valid}), .ready_in_bus({branchC_15_in2_ready, branchC_15_in1_ready}), 
		.data_out_bus({branchC_15_out2_data, branchC_15_out1_data}), .valid_out_bus({branchC_15_out2_valid, branchC_15_out1_valid}), .ready_out_bus({branchC_15_out2_ready, branchC_15_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_0
		(.clk(source_0_clk), .rst(source_0_rst),
		.data_out_bus({source_0_out1_data}), .valid_out_bus({source_0_out1_valid}), .ready_out_bus({source_0_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(5))source_node_source_1
		(.clk(source_1_clk), .rst(source_1_rst),
		.data_out_bus({source_1_out1_data}), .valid_out_bus({source_1_out1_valid}), .ready_out_bus({source_1_out1_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(10), .BB_COUNT(1), .LOAD_COUNT(2), .STORE_COUNT(1))MemCont_MC_A
		(.clk(MC_A_clk), .rst(MC_A_rst),
		.io_storeDataOut(A_dout0), .io_storeAddrOut(A_address0), .io_storeEnable(A_we0),
		.io_loadDataIn(A_din1), .io_loadAddrOut(A_address1), .io_loadEnable(A_ce1),
		.io_bbpValids({MC_A_in1_valid}), .io_bb_stCountArray({MC_A_in1_data}), .io_bbReadyToPrevs({MC_A_in1_ready}), .io_rdPortsPrev_ready({MC_A_in3_ready, MC_A_in2_ready}), .io_rdPortsPrev_valid({MC_A_in3_valid, MC_A_in2_valid}), .io_rdPortsPrev_bits({MC_A_in3_data, MC_A_in2_data}), 	
	.io_wrAddrPorts_ready({MC_A_in4_ready}), .io_wrAddrPorts_valid({MC_A_in4_valid}), .io_wrAddrPorts_bits({MC_A_in4_data}), 	
	.io_wrDataPorts_ready({MC_A_in5_ready}), .io_wrDataPorts_valid({MC_A_in5_valid}), .io_wrDataPorts_bits({MC_A_in5_data}), 	
	.io_rdPortsNext_ready({MC_A_out2_ready, MC_A_out1_ready}), .io_rdPortsNext_valid({MC_A_out2_valid, MC_A_out1_valid}), .io_rdPortsNext_bits({MC_A_out2_data, MC_A_out1_data}), 	
	.io_Empty_Valid({MC_A_out3_valid}), .io_Empty_Ready({MC_A_out3_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(5), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_c
		(.clk(MC_c_clk), .rst(MC_c_rst),
		.io_storeDataOut(c_dout0), .io_storeAddrOut(c_address0), .io_storeEnable(c_we0),
		.io_loadDataIn(c_din1), .io_loadAddrOut(c_address1), .io_loadEnable(c_ce1),
		.io_bbpValids({MC_c_in2_valid}), .io_bb_stCountArray({MC_c_in2_data}), .io_bbReadyToPrevs({MC_c_in2_ready}), .io_rdPortsPrev_ready({MC_c_in1_ready}), .io_rdPortsPrev_valid({MC_c_in1_valid}), .io_rdPortsPrev_bits({MC_c_in1_data}), 	
	.io_wrAddrPorts_ready({MC_c_in3_ready}), .io_wrAddrPorts_valid({MC_c_in3_valid}), .io_wrAddrPorts_bits({MC_c_in3_data}), 	
	.io_wrDataPorts_ready({MC_c_in4_ready}), .io_wrDataPorts_valid({MC_c_in4_valid}), .io_wrDataPorts_bits({MC_c_in4_data}), 	
	.io_rdPortsNext_ready({MC_c_out1_ready}), .io_rdPortsNext_valid({MC_c_out1_valid}), .io_rdPortsNext_bits({MC_c_out1_data}), 	
	.io_Empty_Valid({MC_c_out2_valid}), .io_Empty_Ready({MC_c_out2_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_0
		(.clk(sink_0_clk), .rst(sink_0_rst),
		.data_in_bus({sink_0_in1_data}), .valid_in_bus({sink_0_in1_valid}), .ready_in_bus({sink_0_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_1
		(.clk(sink_1_clk), .rst(sink_1_rst),
		.data_in_bus({sink_1_in1_data}), .valid_in_bus({sink_1_in1_valid}), .ready_in_bus({sink_1_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_2
		(.clk(sink_2_clk), .rst(sink_2_rst),
		.data_in_bus({sink_2_in1_data}), .valid_in_bus({sink_2_in1_valid}), .ready_in_bus({sink_2_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_3
		(.clk(sink_3_clk), .rst(sink_3_rst),
		.data_in_bus({sink_3_in1_data}), .valid_in_bus({sink_3_in1_valid}), .ready_in_bus({sink_3_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_4
		(.clk(sink_4_clk), .rst(sink_4_rst),
		.data_in_bus({sink_4_in1_data}), .valid_in_bus({sink_4_in1_valid}), .ready_in_bus({sink_4_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_5
		(.clk(sink_5_clk), .rst(sink_5_rst),
		.data_in_bus({sink_5_in1_data}), .valid_in_bus({sink_5_in1_valid}), .ready_in_bus({sink_5_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_6
		(.clk(sink_6_clk), .rst(sink_6_rst),
		.data_in_bus({sink_6_in1_data}), .valid_in_bus({sink_6_in1_valid}), .ready_in_bus({sink_6_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_7
		(.clk(sink_7_clk), .rst(sink_7_rst),
		.data_in_bus({sink_7_in1_data}), .valid_in_bus({sink_7_in1_valid}), .ready_in_bus({sink_7_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_8
		(.clk(sink_8_clk), .rst(sink_8_rst),
		.data_in_bus({sink_8_in1_data}), .valid_in_bus({sink_8_in1_valid}), .ready_in_bus({sink_8_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_9
		(.clk(sink_9_clk), .rst(sink_9_rst),
		.data_in_bus({sink_9_in1_data}), .valid_in_bus({sink_9_in1_valid}), .ready_in_bus({sink_9_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_10
		(.clk(sink_10_clk), .rst(sink_10_rst),
		.data_in_bus({sink_10_in1_data}), .valid_in_bus({sink_10_in1_valid}), .ready_in_bus({sink_10_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_11
		(.clk(sink_11_clk), .rst(sink_11_rst),
		.data_in_bus({sink_11_in1_data}), .valid_in_bus({sink_11_in1_valid}), .ready_in_bus({sink_11_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_12
		(.clk(sink_12_clk), .rst(sink_12_rst),
		.data_in_bus({sink_12_in1_data}), .valid_in_bus({sink_12_in1_valid}), .ready_in_bus({sink_12_in1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_100
		(.clk(Buffer_100_clk), .rst(Buffer_100_rst),
		.data_in_bus({Buffer_100_in1_data}), .valid_in_bus({Buffer_100_in1_valid}), .ready_in_bus({Buffer_100_in1_ready}), 
		.data_out_bus({Buffer_100_out1_data}), .valid_out_bus({Buffer_100_out1_valid}), .ready_out_bus({Buffer_100_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_101
		(.clk(Buffer_101_clk), .rst(Buffer_101_rst),
		.data_in_bus({Buffer_101_in1_data}), .valid_in_bus({Buffer_101_in1_valid}), .ready_in_bus({Buffer_101_in1_ready}), 
		.data_out_bus({Buffer_101_out1_data}), .valid_out_bus({Buffer_101_out1_valid}), .ready_out_bus({Buffer_101_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_102
		(.clk(Buffer_102_clk), .rst(Buffer_102_rst),
		.data_in_bus({Buffer_102_in1_data}), .valid_in_bus({Buffer_102_in1_valid}), .ready_in_bus({Buffer_102_in1_ready}), 
		.data_out_bus({Buffer_102_out1_data}), .valid_out_bus({Buffer_102_out1_valid}), .ready_out_bus({Buffer_102_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_103
		(.clk(Buffer_103_clk), .rst(Buffer_103_rst),
		.data_in_bus({Buffer_103_in1_data}), .valid_in_bus({Buffer_103_in1_valid}), .ready_in_bus({Buffer_103_in1_ready}), 
		.data_out_bus({Buffer_103_out1_data}), .valid_out_bus({Buffer_103_out1_valid}), .ready_out_bus({Buffer_103_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_104
		(.clk(Buffer_104_clk), .rst(Buffer_104_rst),
		.data_in_bus({Buffer_104_in1_data}), .valid_in_bus({Buffer_104_in1_valid}), .ready_in_bus({Buffer_104_in1_ready}), 
		.data_out_bus({Buffer_104_out1_data}), .valid_out_bus({Buffer_104_out1_valid}), .ready_out_bus({Buffer_104_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_105
		(.clk(Buffer_105_clk), .rst(Buffer_105_rst),
		.data_in_bus({Buffer_105_in1_data}), .valid_in_bus({Buffer_105_in1_valid}), .ready_in_bus({Buffer_105_in1_ready}), 
		.data_out_bus({Buffer_105_out1_data}), .valid_out_bus({Buffer_105_out1_valid}), .ready_out_bus({Buffer_105_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_106
		(.clk(Buffer_106_clk), .rst(Buffer_106_rst),
		.data_in_bus({Buffer_106_in1_data}), .valid_in_bus({Buffer_106_in1_valid}), .ready_in_bus({Buffer_106_in1_ready}), 
		.data_out_bus({Buffer_106_out1_data}), .valid_out_bus({Buffer_106_out1_valid}), .ready_out_bus({Buffer_106_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_107
		(.clk(Buffer_107_clk), .rst(Buffer_107_rst),
		.data_in_bus({Buffer_107_in1_data}), .valid_in_bus({Buffer_107_in1_valid}), .ready_in_bus({Buffer_107_in1_ready}), 
		.data_out_bus({Buffer_107_out1_data}), .valid_out_bus({Buffer_107_out1_valid}), .ready_out_bus({Buffer_107_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_108
		(.clk(Buffer_108_clk), .rst(Buffer_108_rst),
		.data_in_bus({Buffer_108_in1_data}), .valid_in_bus({Buffer_108_in1_valid}), .ready_in_bus({Buffer_108_in1_ready}), 
		.data_out_bus({Buffer_108_out1_data}), .valid_out_bus({Buffer_108_out1_valid}), .ready_out_bus({Buffer_108_out1_ready}));

endmodule

