module kernel_3mm(
	input clk,
	input rst,

	input [0 : 0]start_in,
	input start_valid,
	output start_ready,

	output [0 : 0]end_out,
	output end_valid,
	input end_ready,

	output [7 : 0]E_address0,
	output E_ce0,
	output E_we0,
	output [31 : 0]E_dout0,
	input [31 : 0]E_din0,
	output [7 : 0]E_address1,
	output E_ce1,
	output E_we1,
	output [31 : 0]E_dout1,
	input [31 : 0]E_din1,

	output [7 : 0]A_address0,
	output A_ce0,
	output A_we0,
	output [31 : 0]A_dout0,
	input [31 : 0]A_din0,
	output [7 : 0]A_address1,
	output A_ce1,
	output A_we1,
	output [31 : 0]A_dout1,
	input [31 : 0]A_din1,

	output [7 : 0]B_address0,
	output B_ce0,
	output B_we0,
	output [31 : 0]B_dout0,
	input [31 : 0]B_din0,
	output [7 : 0]B_address1,
	output B_ce1,
	output B_we1,
	output [31 : 0]B_dout1,
	input [31 : 0]B_din1,

	output [7 : 0]F_address0,
	output F_ce0,
	output F_we0,
	output [31 : 0]F_dout0,
	input [31 : 0]F_din0,
	output [7 : 0]F_address1,
	output F_ce1,
	output F_we1,
	output [31 : 0]F_dout1,
	input [31 : 0]F_din1,

	output [7 : 0]C_address0,
	output C_ce0,
	output C_we0,
	output [31 : 0]C_dout0,
	input [31 : 0]C_din0,
	output [7 : 0]C_address1,
	output C_ce1,
	output C_we1,
	output [31 : 0]C_dout1,
	input [31 : 0]C_din1,

	output [7 : 0]D_address0,
	output D_ce0,
	output D_we0,
	output [31 : 0]D_dout0,
	input [31 : 0]D_din0,
	output [7 : 0]D_address1,
	output D_ce1,
	output D_we1,
	output [31 : 0]D_dout1,
	input [31 : 0]D_din1,

	output [7 : 0]G_address0,
	output G_ce0,
	output G_we0,
	output [31 : 0]G_dout0,
	input [31 : 0]G_din0,
	output [7 : 0]G_address1,
	output G_ce1,
	output G_we1,
	output [31 : 0]G_dout1,
	input [31 : 0]G_din1

);

	wire phi_3_clk;
	wire phi_3_rst;
	wire [0 : 0]phi_3_in1_data;
	wire phi_3_in1_ready;
	wire phi_3_in1_valid;
	wire [3 : 0]phi_3_in2_data;
	wire phi_3_in2_ready;
	wire phi_3_in2_valid;
	wire [3 : 0]phi_3_in3_data;
	wire phi_3_in3_ready;
	wire phi_3_in3_valid;
	wire [3 : 0]phi_3_out1_data;
	wire phi_3_out1_ready;
	wire phi_3_out1_valid;

	wire cst_2_clk;
	wire cst_2_rst;
	wire [1 : 0]cst_2_in1_data;
	wire cst_2_in1_ready;
	wire cst_2_in1_valid;
	wire [1 : 0]cst_2_out1_data;
	wire cst_2_out1_ready;
	wire cst_2_out1_valid;

	wire shl_4_clk;
	wire shl_4_rst;
	wire [6 : 0]shl_4_in1_data;
	wire shl_4_in1_ready;
	wire shl_4_in1_valid;
	wire [6 : 0]shl_4_in2_data;
	wire shl_4_in2_ready;
	wire shl_4_in2_valid;
	wire [6 : 0]shl_4_out1_data;
	wire shl_4_out1_ready;
	wire shl_4_out1_valid;

	wire add_5_clk;
	wire add_5_rst;
	wire [7 : 0]add_5_in1_data;
	wire add_5_in1_ready;
	wire add_5_in1_valid;
	wire [7 : 0]add_5_in2_data;
	wire add_5_in2_ready;
	wire add_5_in2_valid;
	wire [7 : 0]add_5_out1_data;
	wire add_5_out1_ready;
	wire add_5_out1_valid;

	wire load_8_clk;
	wire load_8_rst;
	wire [31 : 0]load_8_in1_data;
	wire load_8_in1_ready;
	wire load_8_in1_valid;
	wire [7 : 0]load_8_in2_data;
	wire load_8_in2_ready;
	wire load_8_in2_valid;
	wire [31 : 0]load_8_out1_data;
	wire load_8_out1_ready;
	wire load_8_out1_valid;
	wire [7 : 0]load_8_out2_data;
	wire load_8_out2_ready;
	wire load_8_out2_valid;

	wire brCst_block3_clk;
	wire brCst_block3_rst;
	wire [0 : 0]brCst_block3_in1_data;
	wire brCst_block3_in1_ready;
	wire brCst_block3_in1_valid;
	wire [0 : 0]brCst_block3_out1_data;
	wire brCst_block3_out1_ready;
	wire brCst_block3_out1_valid;

	wire cst_3_clk;
	wire cst_3_rst;
	wire [0 : 0]cst_3_in1_data;
	wire cst_3_in1_ready;
	wire cst_3_in1_valid;
	wire [0 : 0]cst_3_out1_data;
	wire cst_3_out1_ready;
	wire cst_3_out1_valid;

	wire phi_n4_clk;
	wire phi_n4_rst;
	wire [3 : 0]phi_n4_in1_data;
	wire phi_n4_in1_ready;
	wire phi_n4_in1_valid;
	wire [3 : 0]phi_n4_in2_data;
	wire phi_n4_in2_ready;
	wire phi_n4_in2_valid;
	wire [3 : 0]phi_n4_out1_data;
	wire phi_n4_out1_ready;
	wire phi_n4_out1_valid;

	wire fork_0_clk;
	wire fork_0_rst;
	wire [3 : 0]fork_0_in1_data;
	wire fork_0_in1_ready;
	wire fork_0_in1_valid;
	wire [3 : 0]fork_0_out1_data;
	wire fork_0_out1_ready;
	wire fork_0_out1_valid;
	wire [3 : 0]fork_0_out2_data;
	wire fork_0_out2_ready;
	wire fork_0_out2_valid;

	wire fork_20_clk;
	wire fork_20_rst;
	wire [3 : 0]fork_20_in1_data;
	wire fork_20_in1_ready;
	wire fork_20_in1_valid;
	wire [3 : 0]fork_20_out1_data;
	wire fork_20_out1_ready;
	wire fork_20_out1_valid;
	wire [3 : 0]fork_20_out2_data;
	wire fork_20_out2_ready;
	wire fork_20_out2_valid;

	wire branch_3_clk;
	wire branch_3_rst;
	wire [31 : 0]branch_3_in1_data;
	wire branch_3_in1_ready;
	wire branch_3_in1_valid;
	wire [0 : 0]branch_3_in2_data;
	wire branch_3_in2_ready;
	wire branch_3_in2_valid;
	wire [31 : 0]branch_3_out1_data;
	wire branch_3_out1_ready;
	wire branch_3_out1_valid;
	wire [31 : 0]branch_3_out2_data;
	wire branch_3_out2_ready;
	wire branch_3_out2_valid;

	wire branch_4_clk;
	wire branch_4_rst;
	wire [0 : 0]branch_4_in1_data;
	wire branch_4_in1_ready;
	wire branch_4_in1_valid;
	wire [0 : 0]branch_4_in2_data;
	wire branch_4_in2_ready;
	wire branch_4_in2_valid;
	wire [0 : 0]branch_4_out1_data;
	wire branch_4_out1_ready;
	wire branch_4_out1_valid;
	wire [0 : 0]branch_4_out2_data;
	wire branch_4_out2_ready;
	wire branch_4_out2_valid;

	wire branch_5_clk;
	wire branch_5_rst;
	wire [3 : 0]branch_5_in1_data;
	wire branch_5_in1_ready;
	wire branch_5_in1_valid;
	wire [0 : 0]branch_5_in2_data;
	wire branch_5_in2_ready;
	wire branch_5_in2_valid;
	wire [3 : 0]branch_5_out1_data;
	wire branch_5_out1_ready;
	wire branch_5_out1_valid;
	wire [3 : 0]branch_5_out2_data;
	wire branch_5_out2_ready;
	wire branch_5_out2_valid;

	wire branch_6_clk;
	wire branch_6_rst;
	wire [3 : 0]branch_6_in1_data;
	wire branch_6_in1_ready;
	wire branch_6_in1_valid;
	wire [0 : 0]branch_6_in2_data;
	wire branch_6_in2_ready;
	wire branch_6_in2_valid;
	wire [3 : 0]branch_6_out1_data;
	wire branch_6_out1_ready;
	wire branch_6_out1_valid;
	wire [3 : 0]branch_6_out2_data;
	wire branch_6_out2_ready;
	wire branch_6_out2_valid;

	wire fork_35_clk;
	wire fork_35_rst;
	wire [0 : 0]fork_35_in1_data;
	wire fork_35_in1_ready;
	wire fork_35_in1_valid;
	wire [0 : 0]fork_35_out1_data;
	wire fork_35_out1_ready;
	wire fork_35_out1_valid;
	wire [0 : 0]fork_35_out2_data;
	wire fork_35_out2_ready;
	wire fork_35_out2_valid;
	wire [0 : 0]fork_35_out3_data;
	wire fork_35_out3_ready;
	wire fork_35_out3_valid;
	wire [0 : 0]fork_35_out4_data;
	wire fork_35_out4_ready;
	wire fork_35_out4_valid;
	wire [0 : 0]fork_35_out5_data;
	wire fork_35_out5_ready;
	wire fork_35_out5_valid;

	wire phiC_22_clk;
	wire phiC_22_rst;
	wire [0 : 0]phiC_22_in1_data;
	wire phiC_22_in1_ready;
	wire phiC_22_in1_valid;
	wire [0 : 0]phiC_22_in2_data;
	wire phiC_22_in2_ready;
	wire phiC_22_in2_valid;
	wire [0 : 0]phiC_22_out1_data;
	wire phiC_22_out1_ready;
	wire phiC_22_out1_valid;
	wire [0 : 0]phiC_22_out2_data;
	wire phiC_22_out2_ready;
	wire phiC_22_out2_valid;

	wire forkC_55_clk;
	wire forkC_55_rst;
	wire [0 : 0]forkC_55_in1_data;
	wire forkC_55_in1_ready;
	wire forkC_55_in1_valid;
	wire [0 : 0]forkC_55_out1_data;
	wire forkC_55_out1_ready;
	wire forkC_55_out1_valid;
	wire [0 : 0]forkC_55_out2_data;
	wire forkC_55_out2_ready;
	wire forkC_55_out2_valid;
	wire [0 : 0]forkC_55_out3_data;
	wire forkC_55_out3_ready;
	wire forkC_55_out3_valid;

	wire branchC_44_clk;
	wire branchC_44_rst;
	wire [0 : 0]branchC_44_in1_data;
	wire branchC_44_in1_ready;
	wire branchC_44_in1_valid;
	wire [0 : 0]branchC_44_in2_data;
	wire branchC_44_in2_ready;
	wire branchC_44_in2_valid;
	wire [0 : 0]branchC_44_out1_data;
	wire branchC_44_out1_ready;
	wire branchC_44_out1_valid;
	wire [0 : 0]branchC_44_out2_data;
	wire branchC_44_out2_ready;
	wire branchC_44_out2_valid;

	wire source_0_clk;
	wire source_0_rst;
	wire [1 : 0]source_0_out1_data;
	wire source_0_out1_ready;
	wire source_0_out1_valid;

	wire cst_8_clk;
	wire cst_8_rst;
	wire [1 : 0]cst_8_in1_data;
	wire cst_8_in1_ready;
	wire cst_8_in1_valid;
	wire [1 : 0]cst_8_out1_data;
	wire cst_8_out1_ready;
	wire cst_8_out1_valid;

	wire shl_27_clk;
	wire shl_27_rst;
	wire [6 : 0]shl_27_in1_data;
	wire shl_27_in1_ready;
	wire shl_27_in1_valid;
	wire [6 : 0]shl_27_in2_data;
	wire shl_27_in2_ready;
	wire shl_27_in2_valid;
	wire [6 : 0]shl_27_out1_data;
	wire shl_27_out1_ready;
	wire shl_27_out1_valid;

	wire add_28_clk;
	wire add_28_rst;
	wire [7 : 0]add_28_in1_data;
	wire add_28_in1_ready;
	wire add_28_in1_valid;
	wire [7 : 0]add_28_in2_data;
	wire add_28_in2_ready;
	wire add_28_in2_valid;
	wire [7 : 0]add_28_out1_data;
	wire add_28_out1_ready;
	wire add_28_out1_valid;

	wire store_0_clk;
	wire store_0_rst;
	wire [31 : 0]store_0_in1_data;
	wire store_0_in1_ready;
	wire store_0_in1_valid;
	wire [7 : 0]store_0_in2_data;
	wire store_0_in2_ready;
	wire store_0_in2_valid;
	wire [31 : 0]store_0_out1_data;
	wire store_0_out1_ready;
	wire store_0_out1_valid;
	wire [7 : 0]store_0_out2_data;
	wire store_0_out2_ready;
	wire store_0_out2_valid;

	wire cst_9_clk;
	wire cst_9_rst;
	wire [0 : 0]cst_9_in1_data;
	wire cst_9_in1_ready;
	wire cst_9_in1_valid;
	wire [0 : 0]cst_9_out1_data;
	wire cst_9_out1_ready;
	wire cst_9_out1_valid;

	wire add_31_clk;
	wire add_31_rst;
	wire [3 : 0]add_31_in1_data;
	wire add_31_in1_ready;
	wire add_31_in1_valid;
	wire [3 : 0]add_31_in2_data;
	wire add_31_in2_ready;
	wire add_31_in2_valid;
	wire [3 : 0]add_31_out1_data;
	wire add_31_out1_ready;
	wire add_31_out1_valid;

	wire cst_10_clk;
	wire cst_10_rst;
	wire [3 : 0]cst_10_in1_data;
	wire cst_10_in1_ready;
	wire cst_10_in1_valid;
	wire [3 : 0]cst_10_out1_data;
	wire cst_10_out1_ready;
	wire cst_10_out1_valid;

	wire icmp_32_clk;
	wire icmp_32_rst;
	wire [3 : 0]icmp_32_in1_data;
	wire icmp_32_in1_ready;
	wire icmp_32_in1_valid;
	wire [3 : 0]icmp_32_in2_data;
	wire icmp_32_in2_ready;
	wire icmp_32_in2_valid;
	wire [0 : 0]icmp_32_out1_data;
	wire icmp_32_out1_ready;
	wire icmp_32_out1_valid;

	wire phi_n5_clk;
	wire phi_n5_rst;
	wire [3 : 0]phi_n5_in1_data;
	wire phi_n5_in1_ready;
	wire phi_n5_in1_valid;
	wire [3 : 0]phi_n5_out1_data;
	wire phi_n5_out1_ready;
	wire phi_n5_out1_valid;

	wire phi_n6_clk;
	wire phi_n6_rst;
	wire [3 : 0]phi_n6_in1_data;
	wire phi_n6_in1_ready;
	wire phi_n6_in1_valid;
	wire [3 : 0]phi_n6_out1_data;
	wire phi_n6_out1_ready;
	wire phi_n6_out1_valid;

	wire phi_n7_clk;
	wire phi_n7_rst;
	wire [31 : 0]phi_n7_in1_data;
	wire phi_n7_in1_ready;
	wire phi_n7_in1_valid;
	wire [31 : 0]phi_n7_out1_data;
	wire phi_n7_out1_ready;
	wire phi_n7_out1_valid;

	wire fork_4_clk;
	wire fork_4_rst;
	wire [3 : 0]fork_4_in1_data;
	wire fork_4_in1_ready;
	wire fork_4_in1_valid;
	wire [3 : 0]fork_4_out1_data;
	wire fork_4_out1_ready;
	wire fork_4_out1_valid;
	wire [3 : 0]fork_4_out2_data;
	wire fork_4_out2_ready;
	wire fork_4_out2_valid;

	wire fork_21_clk;
	wire fork_21_rst;
	wire [3 : 0]fork_21_in1_data;
	wire fork_21_in1_ready;
	wire fork_21_in1_valid;
	wire [3 : 0]fork_21_out1_data;
	wire fork_21_out1_ready;
	wire fork_21_out1_valid;
	wire [3 : 0]fork_21_out2_data;
	wire fork_21_out2_ready;
	wire fork_21_out2_valid;

	wire fork_22_clk;
	wire fork_22_rst;
	wire [3 : 0]fork_22_in1_data;
	wire fork_22_in1_ready;
	wire fork_22_in1_valid;
	wire [3 : 0]fork_22_out1_data;
	wire fork_22_out1_ready;
	wire fork_22_out1_valid;
	wire [3 : 0]fork_22_out2_data;
	wire fork_22_out2_ready;
	wire fork_22_out2_valid;

	wire branch_11_clk;
	wire branch_11_rst;
	wire [3 : 0]branch_11_in1_data;
	wire branch_11_in1_ready;
	wire branch_11_in1_valid;
	wire [0 : 0]branch_11_in2_data;
	wire branch_11_in2_ready;
	wire branch_11_in2_valid;
	wire [3 : 0]branch_11_out1_data;
	wire branch_11_out1_ready;
	wire branch_11_out1_valid;
	wire [3 : 0]branch_11_out2_data;
	wire branch_11_out2_ready;
	wire branch_11_out2_valid;

	wire branch_12_clk;
	wire branch_12_rst;
	wire [3 : 0]branch_12_in1_data;
	wire branch_12_in1_ready;
	wire branch_12_in1_valid;
	wire [0 : 0]branch_12_in2_data;
	wire branch_12_in2_ready;
	wire branch_12_in2_valid;
	wire [3 : 0]branch_12_out1_data;
	wire branch_12_out1_ready;
	wire branch_12_out1_valid;
	wire [3 : 0]branch_12_out2_data;
	wire branch_12_out2_ready;
	wire branch_12_out2_valid;

	wire fork_37_clk;
	wire fork_37_rst;
	wire [0 : 0]fork_37_in1_data;
	wire fork_37_in1_ready;
	wire fork_37_in1_valid;
	wire [0 : 0]fork_37_out1_data;
	wire fork_37_out1_ready;
	wire fork_37_out1_valid;
	wire [0 : 0]fork_37_out2_data;
	wire fork_37_out2_ready;
	wire fork_37_out2_valid;
	wire [0 : 0]fork_37_out3_data;
	wire fork_37_out3_ready;
	wire fork_37_out3_valid;

	wire cst_39_clk;
	wire cst_39_rst;
	wire [0 : 0]cst_39_in1_data;
	wire cst_39_in1_ready;
	wire cst_39_in1_valid;
	wire [0 : 0]cst_39_out1_data;
	wire cst_39_out1_ready;
	wire cst_39_out1_valid;

	wire phiC_24_clk;
	wire phiC_24_rst;
	wire [0 : 0]phiC_24_in1_data;
	wire phiC_24_in1_ready;
	wire phiC_24_in1_valid;
	wire [0 : 0]phiC_24_out1_data;
	wire phiC_24_out1_ready;
	wire phiC_24_out1_valid;

	wire forkC_57_clk;
	wire forkC_57_rst;
	wire [0 : 0]forkC_57_in1_data;
	wire forkC_57_in1_ready;
	wire forkC_57_in1_valid;
	wire [0 : 0]forkC_57_out1_data;
	wire forkC_57_out1_ready;
	wire forkC_57_out1_valid;
	wire [0 : 0]forkC_57_out2_data;
	wire forkC_57_out2_ready;
	wire forkC_57_out2_valid;

	wire branchC_46_clk;
	wire branchC_46_rst;
	wire [0 : 0]branchC_46_in1_data;
	wire branchC_46_in1_ready;
	wire branchC_46_in1_valid;
	wire [0 : 0]branchC_46_in2_data;
	wire branchC_46_in2_ready;
	wire branchC_46_in2_valid;
	wire [0 : 0]branchC_46_out1_data;
	wire branchC_46_out1_ready;
	wire branchC_46_out1_valid;
	wire [0 : 0]branchC_46_out2_data;
	wire branchC_46_out2_ready;
	wire branchC_46_out2_valid;

	wire source_5_clk;
	wire source_5_rst;
	wire [1 : 0]source_5_out1_data;
	wire source_5_out1_ready;
	wire source_5_out1_valid;

	wire source_6_clk;
	wire source_6_rst;
	wire [0 : 0]source_6_out1_data;
	wire source_6_out1_ready;
	wire source_6_out1_valid;

	wire source_7_clk;
	wire source_7_rst;
	wire [3 : 0]source_7_out1_data;
	wire source_7_out1_ready;
	wire source_7_out1_valid;

	wire brCst_block1_clk;
	wire brCst_block1_rst;
	wire [0 : 0]brCst_block1_in1_data;
	wire brCst_block1_in1_ready;
	wire brCst_block1_in1_valid;
	wire [0 : 0]brCst_block1_out1_data;
	wire brCst_block1_out1_ready;
	wire brCst_block1_out1_valid;

	wire cst_0_clk;
	wire cst_0_rst;
	wire [0 : 0]cst_0_in1_data;
	wire cst_0_in1_ready;
	wire cst_0_in1_valid;
	wire [0 : 0]cst_0_out1_data;
	wire cst_0_out1_ready;
	wire cst_0_out1_valid;

	wire branch_0_clk;
	wire branch_0_rst;
	wire [0 : 0]branch_0_in1_data;
	wire branch_0_in1_ready;
	wire branch_0_in1_valid;
	wire [0 : 0]branch_0_in2_data;
	wire branch_0_in2_ready;
	wire branch_0_in2_valid;
	wire [0 : 0]branch_0_out1_data;
	wire branch_0_out1_ready;
	wire branch_0_out1_valid;
	wire [0 : 0]branch_0_out2_data;
	wire branch_0_out2_ready;
	wire branch_0_out2_valid;

	wire start_0_clk;
	wire start_0_rst;
	wire [0 : 0]start_0_in1_data;
	wire start_0_in1_ready;
	wire start_0_in1_valid;
	wire [0 : 0]start_0_out1_data;
	wire start_0_out1_ready;
	wire start_0_out1_valid;

	wire forkC_52_clk;
	wire forkC_52_rst;
	wire [0 : 0]forkC_52_in1_data;
	wire forkC_52_in1_ready;
	wire forkC_52_in1_valid;
	wire [0 : 0]forkC_52_out1_data;
	wire forkC_52_out1_ready;
	wire forkC_52_out1_valid;
	wire [0 : 0]forkC_52_out2_data;
	wire forkC_52_out2_ready;
	wire forkC_52_out2_valid;
	wire [0 : 0]forkC_52_out3_data;
	wire forkC_52_out3_ready;
	wire forkC_52_out3_valid;

	wire branchC_42_clk;
	wire branchC_42_rst;
	wire [0 : 0]branchC_42_in1_data;
	wire branchC_42_in1_ready;
	wire branchC_42_in1_valid;
	wire [0 : 0]branchC_42_in2_data;
	wire branchC_42_in2_ready;
	wire branchC_42_in2_valid;
	wire [0 : 0]branchC_42_out1_data;
	wire branchC_42_out1_ready;
	wire branchC_42_out1_valid;
	wire [0 : 0]branchC_42_out2_data;
	wire branchC_42_out2_ready;
	wire branchC_42_out2_valid;

	wire fork_53_clk;
	wire fork_53_rst;
	wire [0 : 0]fork_53_in1_data;
	wire fork_53_in1_ready;
	wire fork_53_in1_valid;
	wire [0 : 0]fork_53_out1_data;
	wire fork_53_out1_ready;
	wire fork_53_out1_valid;
	wire [0 : 0]fork_53_out2_data;
	wire fork_53_out2_ready;
	wire fork_53_out2_valid;

	wire phi_77_clk;
	wire phi_77_rst;
	wire [0 : 0]phi_77_in1_data;
	wire phi_77_in1_ready;
	wire phi_77_in1_valid;
	wire [3 : 0]phi_77_in2_data;
	wire phi_77_in2_ready;
	wire phi_77_in2_valid;
	wire [3 : 0]phi_77_in3_data;
	wire phi_77_in3_ready;
	wire phi_77_in3_valid;
	wire [3 : 0]phi_77_out1_data;
	wire phi_77_out1_ready;
	wire phi_77_out1_valid;

	wire cst_28_clk;
	wire cst_28_rst;
	wire [1 : 0]cst_28_in1_data;
	wire cst_28_in1_ready;
	wire cst_28_in1_valid;
	wire [1 : 0]cst_28_out1_data;
	wire cst_28_out1_ready;
	wire cst_28_out1_valid;

	wire shl_78_clk;
	wire shl_78_rst;
	wire [6 : 0]shl_78_in1_data;
	wire shl_78_in1_ready;
	wire shl_78_in1_valid;
	wire [6 : 0]shl_78_in2_data;
	wire shl_78_in2_ready;
	wire shl_78_in2_valid;
	wire [6 : 0]shl_78_out1_data;
	wire shl_78_out1_ready;
	wire shl_78_out1_valid;

	wire add_79_clk;
	wire add_79_rst;
	wire [7 : 0]add_79_in1_data;
	wire add_79_in1_ready;
	wire add_79_in1_valid;
	wire [7 : 0]add_79_in2_data;
	wire add_79_in2_ready;
	wire add_79_in2_valid;
	wire [7 : 0]add_79_out1_data;
	wire add_79_out1_ready;
	wire add_79_out1_valid;

	wire load_82_clk;
	wire load_82_rst;
	wire [31 : 0]load_82_in1_data;
	wire load_82_in1_ready;
	wire load_82_in1_valid;
	wire [7 : 0]load_82_in2_data;
	wire load_82_in2_ready;
	wire load_82_in2_valid;
	wire [31 : 0]load_82_out1_data;
	wire load_82_out1_ready;
	wire load_82_out1_valid;
	wire [7 : 0]load_82_out2_data;
	wire load_82_out2_ready;
	wire load_82_out2_valid;

	wire brCst_block15_clk;
	wire brCst_block15_rst;
	wire [0 : 0]brCst_block15_in1_data;
	wire brCst_block15_in1_ready;
	wire brCst_block15_in1_valid;
	wire [0 : 0]brCst_block15_out1_data;
	wire brCst_block15_out1_ready;
	wire brCst_block15_out1_valid;

	wire cst_29_clk;
	wire cst_29_rst;
	wire [0 : 0]cst_29_in1_data;
	wire cst_29_in1_ready;
	wire cst_29_in1_valid;
	wire [0 : 0]cst_29_out1_data;
	wire cst_29_out1_ready;
	wire cst_29_out1_valid;

	wire phi_n15_clk;
	wire phi_n15_rst;
	wire [3 : 0]phi_n15_in1_data;
	wire phi_n15_in1_ready;
	wire phi_n15_in1_valid;
	wire [3 : 0]phi_n15_in2_data;
	wire phi_n15_in2_ready;
	wire phi_n15_in2_valid;
	wire [3 : 0]phi_n15_out1_data;
	wire phi_n15_out1_ready;
	wire phi_n15_out1_valid;

	wire fork_12_clk;
	wire fork_12_rst;
	wire [3 : 0]fork_12_in1_data;
	wire fork_12_in1_ready;
	wire fork_12_in1_valid;
	wire [3 : 0]fork_12_out1_data;
	wire fork_12_out1_ready;
	wire fork_12_out1_valid;
	wire [3 : 0]fork_12_out2_data;
	wire fork_12_out2_ready;
	wire fork_12_out2_valid;

	wire fork_28_clk;
	wire fork_28_rst;
	wire [3 : 0]fork_28_in1_data;
	wire fork_28_in1_ready;
	wire fork_28_in1_valid;
	wire [3 : 0]fork_28_out1_data;
	wire fork_28_out1_ready;
	wire fork_28_out1_valid;
	wire [3 : 0]fork_28_out2_data;
	wire fork_28_out2_ready;
	wire fork_28_out2_valid;

	wire branch_31_clk;
	wire branch_31_rst;
	wire [31 : 0]branch_31_in1_data;
	wire branch_31_in1_ready;
	wire branch_31_in1_valid;
	wire [0 : 0]branch_31_in2_data;
	wire branch_31_in2_ready;
	wire branch_31_in2_valid;
	wire [31 : 0]branch_31_out1_data;
	wire branch_31_out1_ready;
	wire branch_31_out1_valid;
	wire [31 : 0]branch_31_out2_data;
	wire branch_31_out2_ready;
	wire branch_31_out2_valid;

	wire branch_32_clk;
	wire branch_32_rst;
	wire [0 : 0]branch_32_in1_data;
	wire branch_32_in1_ready;
	wire branch_32_in1_valid;
	wire [0 : 0]branch_32_in2_data;
	wire branch_32_in2_ready;
	wire branch_32_in2_valid;
	wire [0 : 0]branch_32_out1_data;
	wire branch_32_out1_ready;
	wire branch_32_out1_valid;
	wire [0 : 0]branch_32_out2_data;
	wire branch_32_out2_ready;
	wire branch_32_out2_valid;

	wire branch_33_clk;
	wire branch_33_rst;
	wire [3 : 0]branch_33_in1_data;
	wire branch_33_in1_ready;
	wire branch_33_in1_valid;
	wire [0 : 0]branch_33_in2_data;
	wire branch_33_in2_ready;
	wire branch_33_in2_valid;
	wire [3 : 0]branch_33_out1_data;
	wire branch_33_out1_ready;
	wire branch_33_out1_valid;
	wire [3 : 0]branch_33_out2_data;
	wire branch_33_out2_ready;
	wire branch_33_out2_valid;

	wire branch_34_clk;
	wire branch_34_rst;
	wire [3 : 0]branch_34_in1_data;
	wire branch_34_in1_ready;
	wire branch_34_in1_valid;
	wire [0 : 0]branch_34_in2_data;
	wire branch_34_in2_ready;
	wire branch_34_in2_valid;
	wire [3 : 0]branch_34_out1_data;
	wire branch_34_out1_ready;
	wire branch_34_out1_valid;
	wire [3 : 0]branch_34_out2_data;
	wire branch_34_out2_ready;
	wire branch_34_out2_valid;

	wire fork_47_clk;
	wire fork_47_rst;
	wire [0 : 0]fork_47_in1_data;
	wire fork_47_in1_ready;
	wire fork_47_in1_valid;
	wire [0 : 0]fork_47_out1_data;
	wire fork_47_out1_ready;
	wire fork_47_out1_valid;
	wire [0 : 0]fork_47_out2_data;
	wire fork_47_out2_ready;
	wire fork_47_out2_valid;
	wire [0 : 0]fork_47_out3_data;
	wire fork_47_out3_ready;
	wire fork_47_out3_valid;
	wire [0 : 0]fork_47_out4_data;
	wire fork_47_out4_ready;
	wire fork_47_out4_valid;
	wire [0 : 0]fork_47_out5_data;
	wire fork_47_out5_ready;
	wire fork_47_out5_valid;

	wire phiC_34_clk;
	wire phiC_34_rst;
	wire [0 : 0]phiC_34_in1_data;
	wire phiC_34_in1_ready;
	wire phiC_34_in1_valid;
	wire [0 : 0]phiC_34_in2_data;
	wire phiC_34_in2_ready;
	wire phiC_34_in2_valid;
	wire [0 : 0]phiC_34_out1_data;
	wire phiC_34_out1_ready;
	wire phiC_34_out1_valid;
	wire [0 : 0]phiC_34_out2_data;
	wire phiC_34_out2_ready;
	wire phiC_34_out2_valid;

	wire forkC_71_clk;
	wire forkC_71_rst;
	wire [0 : 0]forkC_71_in1_data;
	wire forkC_71_in1_ready;
	wire forkC_71_in1_valid;
	wire [0 : 0]forkC_71_out1_data;
	wire forkC_71_out1_ready;
	wire forkC_71_out1_valid;
	wire [0 : 0]forkC_71_out2_data;
	wire forkC_71_out2_ready;
	wire forkC_71_out2_valid;
	wire [0 : 0]forkC_71_out3_data;
	wire forkC_71_out3_ready;
	wire forkC_71_out3_valid;

	wire branchC_56_clk;
	wire branchC_56_rst;
	wire [0 : 0]branchC_56_in1_data;
	wire branchC_56_in1_ready;
	wire branchC_56_in1_valid;
	wire [0 : 0]branchC_56_in2_data;
	wire branchC_56_in2_ready;
	wire branchC_56_in2_valid;
	wire [0 : 0]branchC_56_out1_data;
	wire branchC_56_out1_ready;
	wire branchC_56_out1_valid;
	wire [0 : 0]branchC_56_out2_data;
	wire branchC_56_out2_ready;
	wire branchC_56_out2_valid;

	wire source_20_clk;
	wire source_20_rst;
	wire [1 : 0]source_20_out1_data;
	wire source_20_out1_ready;
	wire source_20_out1_valid;

	wire phi_38_clk;
	wire phi_38_rst;
	wire [0 : 0]phi_38_in1_data;
	wire phi_38_in1_ready;
	wire phi_38_in1_valid;
	wire [3 : 0]phi_38_in2_data;
	wire phi_38_in2_ready;
	wire phi_38_in2_valid;
	wire [3 : 0]phi_38_in3_data;
	wire phi_38_in3_ready;
	wire phi_38_in3_valid;
	wire [3 : 0]phi_38_out1_data;
	wire phi_38_out1_ready;
	wire phi_38_out1_valid;

	wire brCst_block8_clk;
	wire brCst_block8_rst;
	wire [0 : 0]brCst_block8_in1_data;
	wire brCst_block8_in1_ready;
	wire brCst_block8_in1_valid;
	wire [0 : 0]brCst_block8_out1_data;
	wire brCst_block8_out1_ready;
	wire brCst_block8_out1_valid;

	wire cst_14_clk;
	wire cst_14_rst;
	wire [0 : 0]cst_14_in1_data;
	wire cst_14_in1_ready;
	wire cst_14_in1_valid;
	wire [0 : 0]cst_14_out1_data;
	wire cst_14_out1_ready;
	wire cst_14_out1_valid;

	wire branch_15_clk;
	wire branch_15_rst;
	wire [0 : 0]branch_15_in1_data;
	wire branch_15_in1_ready;
	wire branch_15_in1_valid;
	wire [0 : 0]branch_15_in2_data;
	wire branch_15_in2_ready;
	wire branch_15_in2_valid;
	wire [0 : 0]branch_15_out1_data;
	wire branch_15_out1_ready;
	wire branch_15_out1_valid;
	wire [0 : 0]branch_15_out2_data;
	wire branch_15_out2_ready;
	wire branch_15_out2_valid;

	wire branch_16_clk;
	wire branch_16_rst;
	wire [3 : 0]branch_16_in1_data;
	wire branch_16_in1_ready;
	wire branch_16_in1_valid;
	wire [0 : 0]branch_16_in2_data;
	wire branch_16_in2_ready;
	wire branch_16_in2_valid;
	wire [3 : 0]branch_16_out1_data;
	wire branch_16_out1_ready;
	wire branch_16_out1_valid;
	wire [3 : 0]branch_16_out2_data;
	wire branch_16_out2_ready;
	wire branch_16_out2_valid;

	wire fork_40_clk;
	wire fork_40_rst;
	wire [0 : 0]fork_40_in1_data;
	wire fork_40_in1_ready;
	wire fork_40_in1_valid;
	wire [0 : 0]fork_40_out1_data;
	wire fork_40_out1_ready;
	wire fork_40_out1_valid;
	wire [0 : 0]fork_40_out2_data;
	wire fork_40_out2_ready;
	wire fork_40_out2_valid;
	wire [0 : 0]fork_40_out3_data;
	wire fork_40_out3_ready;
	wire fork_40_out3_valid;

	wire phiC_27_clk;
	wire phiC_27_rst;
	wire [0 : 0]phiC_27_in1_data;
	wire phiC_27_in1_ready;
	wire phiC_27_in1_valid;
	wire [0 : 0]phiC_27_in2_data;
	wire phiC_27_in2_ready;
	wire phiC_27_in2_valid;
	wire [0 : 0]phiC_27_out1_data;
	wire phiC_27_out1_ready;
	wire phiC_27_out1_valid;
	wire [0 : 0]phiC_27_out2_data;
	wire phiC_27_out2_ready;
	wire phiC_27_out2_valid;

	wire forkC_62_clk;
	wire forkC_62_rst;
	wire [0 : 0]forkC_62_in1_data;
	wire forkC_62_in1_ready;
	wire forkC_62_in1_valid;
	wire [0 : 0]forkC_62_out1_data;
	wire forkC_62_out1_ready;
	wire forkC_62_out1_valid;
	wire [0 : 0]forkC_62_out2_data;
	wire forkC_62_out2_ready;
	wire forkC_62_out2_valid;
	wire [0 : 0]forkC_62_out3_data;
	wire forkC_62_out3_ready;
	wire forkC_62_out3_valid;

	wire branchC_49_clk;
	wire branchC_49_rst;
	wire [0 : 0]branchC_49_in1_data;
	wire branchC_49_in1_ready;
	wire branchC_49_in1_valid;
	wire [0 : 0]branchC_49_in2_data;
	wire branchC_49_in2_ready;
	wire branchC_49_in2_valid;
	wire [0 : 0]branchC_49_out1_data;
	wire branchC_49_out1_ready;
	wire branchC_49_out1_valid;
	wire [0 : 0]branchC_49_out2_data;
	wire branchC_49_out2_ready;
	wire branchC_49_out2_valid;

	wire cst_11_clk;
	wire cst_11_rst;
	wire [0 : 0]cst_11_in1_data;
	wire cst_11_in1_ready;
	wire cst_11_in1_valid;
	wire [0 : 0]cst_11_out1_data;
	wire cst_11_out1_ready;
	wire cst_11_out1_valid;

	wire add_34_clk;
	wire add_34_rst;
	wire [3 : 0]add_34_in1_data;
	wire add_34_in1_ready;
	wire add_34_in1_valid;
	wire [3 : 0]add_34_in2_data;
	wire add_34_in2_ready;
	wire add_34_in2_valid;
	wire [3 : 0]add_34_out1_data;
	wire add_34_out1_ready;
	wire add_34_out1_valid;

	wire cst_12_clk;
	wire cst_12_rst;
	wire [3 : 0]cst_12_in1_data;
	wire cst_12_in1_ready;
	wire cst_12_in1_valid;
	wire [3 : 0]cst_12_out1_data;
	wire cst_12_out1_ready;
	wire cst_12_out1_valid;

	wire icmp_35_clk;
	wire icmp_35_rst;
	wire [3 : 0]icmp_35_in1_data;
	wire icmp_35_in1_ready;
	wire icmp_35_in1_valid;
	wire [3 : 0]icmp_35_in2_data;
	wire icmp_35_in2_ready;
	wire icmp_35_in2_valid;
	wire [0 : 0]icmp_35_out1_data;
	wire icmp_35_out1_ready;
	wire icmp_35_out1_valid;

	wire phi_n3_clk;
	wire phi_n3_rst;
	wire [3 : 0]phi_n3_in1_data;
	wire phi_n3_in1_ready;
	wire phi_n3_in1_valid;
	wire [3 : 0]phi_n3_out1_data;
	wire phi_n3_out1_ready;
	wire phi_n3_out1_valid;

	wire fork_5_clk;
	wire fork_5_rst;
	wire [3 : 0]fork_5_in1_data;
	wire fork_5_in1_ready;
	wire fork_5_in1_valid;
	wire [3 : 0]fork_5_out1_data;
	wire fork_5_out1_ready;
	wire fork_5_out1_valid;
	wire [3 : 0]fork_5_out2_data;
	wire fork_5_out2_ready;
	wire fork_5_out2_valid;

	wire branch_13_clk;
	wire branch_13_rst;
	wire [3 : 0]branch_13_in1_data;
	wire branch_13_in1_ready;
	wire branch_13_in1_valid;
	wire [0 : 0]branch_13_in2_data;
	wire branch_13_in2_ready;
	wire branch_13_in2_valid;
	wire [3 : 0]branch_13_out1_data;
	wire branch_13_out1_ready;
	wire branch_13_out1_valid;
	wire [3 : 0]branch_13_out2_data;
	wire branch_13_out2_ready;
	wire branch_13_out2_valid;

	wire phiC_25_clk;
	wire phiC_25_rst;
	wire [0 : 0]phiC_25_in1_data;
	wire phiC_25_in1_ready;
	wire phiC_25_in1_valid;
	wire [0 : 0]phiC_25_out1_data;
	wire phiC_25_out1_ready;
	wire phiC_25_out1_valid;

	wire branchC_47_clk;
	wire branchC_47_rst;
	wire [0 : 0]branchC_47_in1_data;
	wire branchC_47_in1_ready;
	wire branchC_47_in1_valid;
	wire [0 : 0]branchC_47_in2_data;
	wire branchC_47_in2_ready;
	wire branchC_47_in2_valid;
	wire [0 : 0]branchC_47_out1_data;
	wire branchC_47_out1_ready;
	wire branchC_47_out1_valid;
	wire [0 : 0]branchC_47_out2_data;
	wire branchC_47_out2_ready;
	wire branchC_47_out2_valid;

	wire fork_59_clk;
	wire fork_59_rst;
	wire [0 : 0]fork_59_in1_data;
	wire fork_59_in1_ready;
	wire fork_59_in1_valid;
	wire [0 : 0]fork_59_out1_data;
	wire fork_59_out1_ready;
	wire fork_59_out1_valid;
	wire [0 : 0]fork_59_out2_data;
	wire fork_59_out2_ready;
	wire fork_59_out2_valid;

	wire source_8_clk;
	wire source_8_rst;
	wire [0 : 0]source_8_out1_data;
	wire source_8_out1_ready;
	wire source_8_out1_valid;

	wire source_9_clk;
	wire source_9_rst;
	wire [3 : 0]source_9_out1_data;
	wire source_9_out1_ready;
	wire source_9_out1_valid;

	wire cst_34_clk;
	wire cst_34_rst;
	wire [1 : 0]cst_34_in1_data;
	wire cst_34_in1_ready;
	wire cst_34_in1_valid;
	wire [1 : 0]cst_34_out1_data;
	wire cst_34_out1_ready;
	wire cst_34_out1_valid;

	wire shl_101_clk;
	wire shl_101_rst;
	wire [6 : 0]shl_101_in1_data;
	wire shl_101_in1_ready;
	wire shl_101_in1_valid;
	wire [6 : 0]shl_101_in2_data;
	wire shl_101_in2_ready;
	wire shl_101_in2_valid;
	wire [6 : 0]shl_101_out1_data;
	wire shl_101_out1_ready;
	wire shl_101_out1_valid;

	wire add_102_clk;
	wire add_102_rst;
	wire [7 : 0]add_102_in1_data;
	wire add_102_in1_ready;
	wire add_102_in1_valid;
	wire [7 : 0]add_102_in2_data;
	wire add_102_in2_ready;
	wire add_102_in2_valid;
	wire [7 : 0]add_102_out1_data;
	wire add_102_out1_ready;
	wire add_102_out1_valid;

	wire store_2_clk;
	wire store_2_rst;
	wire [31 : 0]store_2_in1_data;
	wire store_2_in1_ready;
	wire store_2_in1_valid;
	wire [7 : 0]store_2_in2_data;
	wire store_2_in2_ready;
	wire store_2_in2_valid;
	wire [31 : 0]store_2_out1_data;
	wire store_2_out1_ready;
	wire store_2_out1_valid;
	wire [7 : 0]store_2_out2_data;
	wire store_2_out2_ready;
	wire store_2_out2_valid;

	wire cst_35_clk;
	wire cst_35_rst;
	wire [0 : 0]cst_35_in1_data;
	wire cst_35_in1_ready;
	wire cst_35_in1_valid;
	wire [0 : 0]cst_35_out1_data;
	wire cst_35_out1_ready;
	wire cst_35_out1_valid;

	wire add_105_clk;
	wire add_105_rst;
	wire [3 : 0]add_105_in1_data;
	wire add_105_in1_ready;
	wire add_105_in1_valid;
	wire [3 : 0]add_105_in2_data;
	wire add_105_in2_ready;
	wire add_105_in2_valid;
	wire [3 : 0]add_105_out1_data;
	wire add_105_out1_ready;
	wire add_105_out1_valid;

	wire cst_36_clk;
	wire cst_36_rst;
	wire [3 : 0]cst_36_in1_data;
	wire cst_36_in1_ready;
	wire cst_36_in1_valid;
	wire [3 : 0]cst_36_out1_data;
	wire cst_36_out1_ready;
	wire cst_36_out1_valid;

	wire icmp_106_clk;
	wire icmp_106_rst;
	wire [3 : 0]icmp_106_in1_data;
	wire icmp_106_in1_ready;
	wire icmp_106_in1_valid;
	wire [3 : 0]icmp_106_in2_data;
	wire icmp_106_in2_ready;
	wire icmp_106_in2_valid;
	wire [0 : 0]icmp_106_out1_data;
	wire icmp_106_out1_ready;
	wire icmp_106_out1_valid;

	wire phi_n16_clk;
	wire phi_n16_rst;
	wire [3 : 0]phi_n16_in1_data;
	wire phi_n16_in1_ready;
	wire phi_n16_in1_valid;
	wire [3 : 0]phi_n16_out1_data;
	wire phi_n16_out1_ready;
	wire phi_n16_out1_valid;

	wire phi_n17_clk;
	wire phi_n17_rst;
	wire [3 : 0]phi_n17_in1_data;
	wire phi_n17_in1_ready;
	wire phi_n17_in1_valid;
	wire [3 : 0]phi_n17_out1_data;
	wire phi_n17_out1_ready;
	wire phi_n17_out1_valid;

	wire phi_n18_clk;
	wire phi_n18_rst;
	wire [31 : 0]phi_n18_in1_data;
	wire phi_n18_in1_ready;
	wire phi_n18_in1_valid;
	wire [31 : 0]phi_n18_out1_data;
	wire phi_n18_out1_ready;
	wire phi_n18_out1_valid;

	wire fork_16_clk;
	wire fork_16_rst;
	wire [3 : 0]fork_16_in1_data;
	wire fork_16_in1_ready;
	wire fork_16_in1_valid;
	wire [3 : 0]fork_16_out1_data;
	wire fork_16_out1_ready;
	wire fork_16_out1_valid;
	wire [3 : 0]fork_16_out2_data;
	wire fork_16_out2_ready;
	wire fork_16_out2_valid;

	wire fork_29_clk;
	wire fork_29_rst;
	wire [3 : 0]fork_29_in1_data;
	wire fork_29_in1_ready;
	wire fork_29_in1_valid;
	wire [3 : 0]fork_29_out1_data;
	wire fork_29_out1_ready;
	wire fork_29_out1_valid;
	wire [3 : 0]fork_29_out2_data;
	wire fork_29_out2_ready;
	wire fork_29_out2_valid;

	wire fork_30_clk;
	wire fork_30_rst;
	wire [3 : 0]fork_30_in1_data;
	wire fork_30_in1_ready;
	wire fork_30_in1_valid;
	wire [3 : 0]fork_30_out1_data;
	wire fork_30_out1_ready;
	wire fork_30_out1_valid;
	wire [3 : 0]fork_30_out2_data;
	wire fork_30_out2_ready;
	wire fork_30_out2_valid;

	wire branch_39_clk;
	wire branch_39_rst;
	wire [3 : 0]branch_39_in1_data;
	wire branch_39_in1_ready;
	wire branch_39_in1_valid;
	wire [0 : 0]branch_39_in2_data;
	wire branch_39_in2_ready;
	wire branch_39_in2_valid;
	wire [3 : 0]branch_39_out1_data;
	wire branch_39_out1_ready;
	wire branch_39_out1_valid;
	wire [3 : 0]branch_39_out2_data;
	wire branch_39_out2_ready;
	wire branch_39_out2_valid;

	wire branch_40_clk;
	wire branch_40_rst;
	wire [3 : 0]branch_40_in1_data;
	wire branch_40_in1_ready;
	wire branch_40_in1_valid;
	wire [0 : 0]branch_40_in2_data;
	wire branch_40_in2_ready;
	wire branch_40_in2_valid;
	wire [3 : 0]branch_40_out1_data;
	wire branch_40_out1_ready;
	wire branch_40_out1_valid;
	wire [3 : 0]branch_40_out2_data;
	wire branch_40_out2_ready;
	wire branch_40_out2_valid;

	wire fork_49_clk;
	wire fork_49_rst;
	wire [0 : 0]fork_49_in1_data;
	wire fork_49_in1_ready;
	wire fork_49_in1_valid;
	wire [0 : 0]fork_49_out1_data;
	wire fork_49_out1_ready;
	wire fork_49_out1_valid;
	wire [0 : 0]fork_49_out2_data;
	wire fork_49_out2_ready;
	wire fork_49_out2_valid;
	wire [0 : 0]fork_49_out3_data;
	wire fork_49_out3_ready;
	wire fork_49_out3_valid;

	wire cst_41_clk;
	wire cst_41_rst;
	wire [0 : 0]cst_41_in1_data;
	wire cst_41_in1_ready;
	wire cst_41_in1_valid;
	wire [0 : 0]cst_41_out1_data;
	wire cst_41_out1_ready;
	wire cst_41_out1_valid;

	wire phiC_36_clk;
	wire phiC_36_rst;
	wire [0 : 0]phiC_36_in1_data;
	wire phiC_36_in1_ready;
	wire phiC_36_in1_valid;
	wire [0 : 0]phiC_36_out1_data;
	wire phiC_36_out1_ready;
	wire phiC_36_out1_valid;

	wire forkC_73_clk;
	wire forkC_73_rst;
	wire [0 : 0]forkC_73_in1_data;
	wire forkC_73_in1_ready;
	wire forkC_73_in1_valid;
	wire [0 : 0]forkC_73_out1_data;
	wire forkC_73_out1_ready;
	wire forkC_73_out1_valid;
	wire [0 : 0]forkC_73_out2_data;
	wire forkC_73_out2_ready;
	wire forkC_73_out2_valid;

	wire branchC_58_clk;
	wire branchC_58_rst;
	wire [0 : 0]branchC_58_in1_data;
	wire branchC_58_in1_ready;
	wire branchC_58_in1_valid;
	wire [0 : 0]branchC_58_in2_data;
	wire branchC_58_in2_ready;
	wire branchC_58_in2_valid;
	wire [0 : 0]branchC_58_out1_data;
	wire branchC_58_out1_ready;
	wire branchC_58_out1_valid;
	wire [0 : 0]branchC_58_out2_data;
	wire branchC_58_out2_ready;
	wire branchC_58_out2_valid;

	wire source_25_clk;
	wire source_25_rst;
	wire [1 : 0]source_25_out1_data;
	wire source_25_out1_ready;
	wire source_25_out1_valid;

	wire source_26_clk;
	wire source_26_rst;
	wire [0 : 0]source_26_out1_data;
	wire source_26_out1_ready;
	wire source_26_out1_valid;

	wire source_27_clk;
	wire source_27_rst;
	wire [3 : 0]source_27_out1_data;
	wire source_27_out1_ready;
	wire source_27_out1_valid;

	wire cst_21_clk;
	wire cst_21_rst;
	wire [1 : 0]cst_21_in1_data;
	wire cst_21_in1_ready;
	wire cst_21_in1_valid;
	wire [1 : 0]cst_21_out1_data;
	wire cst_21_out1_ready;
	wire cst_21_out1_valid;

	wire shl_64_clk;
	wire shl_64_rst;
	wire [6 : 0]shl_64_in1_data;
	wire shl_64_in1_ready;
	wire shl_64_in1_valid;
	wire [6 : 0]shl_64_in2_data;
	wire shl_64_in2_ready;
	wire shl_64_in2_valid;
	wire [6 : 0]shl_64_out1_data;
	wire shl_64_out1_ready;
	wire shl_64_out1_valid;

	wire add_65_clk;
	wire add_65_rst;
	wire [7 : 0]add_65_in1_data;
	wire add_65_in1_ready;
	wire add_65_in1_valid;
	wire [7 : 0]add_65_in2_data;
	wire add_65_in2_ready;
	wire add_65_in2_valid;
	wire [7 : 0]add_65_out1_data;
	wire add_65_out1_ready;
	wire add_65_out1_valid;

	wire store_1_clk;
	wire store_1_rst;
	wire [31 : 0]store_1_in1_data;
	wire store_1_in1_ready;
	wire store_1_in1_valid;
	wire [7 : 0]store_1_in2_data;
	wire store_1_in2_ready;
	wire store_1_in2_valid;
	wire [31 : 0]store_1_out1_data;
	wire store_1_out1_ready;
	wire store_1_out1_valid;
	wire [7 : 0]store_1_out2_data;
	wire store_1_out2_ready;
	wire store_1_out2_valid;

	wire cst_22_clk;
	wire cst_22_rst;
	wire [0 : 0]cst_22_in1_data;
	wire cst_22_in1_ready;
	wire cst_22_in1_valid;
	wire [0 : 0]cst_22_out1_data;
	wire cst_22_out1_ready;
	wire cst_22_out1_valid;

	wire add_68_clk;
	wire add_68_rst;
	wire [3 : 0]add_68_in1_data;
	wire add_68_in1_ready;
	wire add_68_in1_valid;
	wire [3 : 0]add_68_in2_data;
	wire add_68_in2_ready;
	wire add_68_in2_valid;
	wire [3 : 0]add_68_out1_data;
	wire add_68_out1_ready;
	wire add_68_out1_valid;

	wire cst_23_clk;
	wire cst_23_rst;
	wire [3 : 0]cst_23_in1_data;
	wire cst_23_in1_ready;
	wire cst_23_in1_valid;
	wire [3 : 0]cst_23_out1_data;
	wire cst_23_out1_ready;
	wire cst_23_out1_valid;

	wire icmp_69_clk;
	wire icmp_69_rst;
	wire [3 : 0]icmp_69_in1_data;
	wire icmp_69_in1_ready;
	wire icmp_69_in1_valid;
	wire [3 : 0]icmp_69_in2_data;
	wire icmp_69_in2_ready;
	wire icmp_69_in2_valid;
	wire [0 : 0]icmp_69_out1_data;
	wire icmp_69_out1_ready;
	wire icmp_69_out1_valid;

	wire phi_n0_clk;
	wire phi_n0_rst;
	wire [3 : 0]phi_n0_in1_data;
	wire phi_n0_in1_ready;
	wire phi_n0_in1_valid;
	wire [3 : 0]phi_n0_out1_data;
	wire phi_n0_out1_ready;
	wire phi_n0_out1_valid;

	wire phi_n1_clk;
	wire phi_n1_rst;
	wire [3 : 0]phi_n1_in1_data;
	wire phi_n1_in1_ready;
	wire phi_n1_in1_valid;
	wire [3 : 0]phi_n1_out1_data;
	wire phi_n1_out1_ready;
	wire phi_n1_out1_valid;

	wire phi_n2_clk;
	wire phi_n2_rst;
	wire [31 : 0]phi_n2_in1_data;
	wire phi_n2_in1_ready;
	wire phi_n2_in1_valid;
	wire [31 : 0]phi_n2_out1_data;
	wire phi_n2_out1_ready;
	wire phi_n2_out1_valid;

	wire fork_10_clk;
	wire fork_10_rst;
	wire [3 : 0]fork_10_in1_data;
	wire fork_10_in1_ready;
	wire fork_10_in1_valid;
	wire [3 : 0]fork_10_out1_data;
	wire fork_10_out1_ready;
	wire fork_10_out1_valid;
	wire [3 : 0]fork_10_out2_data;
	wire fork_10_out2_ready;
	wire fork_10_out2_valid;

	wire fork_18_clk;
	wire fork_18_rst;
	wire [3 : 0]fork_18_in1_data;
	wire fork_18_in1_ready;
	wire fork_18_in1_valid;
	wire [3 : 0]fork_18_out1_data;
	wire fork_18_out1_ready;
	wire fork_18_out1_valid;
	wire [3 : 0]fork_18_out2_data;
	wire fork_18_out2_ready;
	wire fork_18_out2_valid;

	wire fork_19_clk;
	wire fork_19_rst;
	wire [3 : 0]fork_19_in1_data;
	wire fork_19_in1_ready;
	wire fork_19_in1_valid;
	wire [3 : 0]fork_19_out1_data;
	wire fork_19_out1_ready;
	wire fork_19_out1_valid;
	wire [3 : 0]fork_19_out2_data;
	wire fork_19_out2_ready;
	wire fork_19_out2_valid;

	wire branch_25_clk;
	wire branch_25_rst;
	wire [3 : 0]branch_25_in1_data;
	wire branch_25_in1_ready;
	wire branch_25_in1_valid;
	wire [0 : 0]branch_25_in2_data;
	wire branch_25_in2_ready;
	wire branch_25_in2_valid;
	wire [3 : 0]branch_25_out1_data;
	wire branch_25_out1_ready;
	wire branch_25_out1_valid;
	wire [3 : 0]branch_25_out2_data;
	wire branch_25_out2_ready;
	wire branch_25_out2_valid;

	wire branch_26_clk;
	wire branch_26_rst;
	wire [3 : 0]branch_26_in1_data;
	wire branch_26_in1_ready;
	wire branch_26_in1_valid;
	wire [0 : 0]branch_26_in2_data;
	wire branch_26_in2_ready;
	wire branch_26_in2_valid;
	wire [3 : 0]branch_26_out1_data;
	wire branch_26_out1_ready;
	wire branch_26_out1_valid;
	wire [3 : 0]branch_26_out2_data;
	wire branch_26_out2_ready;
	wire branch_26_out2_valid;

	wire fork_43_clk;
	wire fork_43_rst;
	wire [0 : 0]fork_43_in1_data;
	wire fork_43_in1_ready;
	wire fork_43_in1_valid;
	wire [0 : 0]fork_43_out1_data;
	wire fork_43_out1_ready;
	wire fork_43_out1_valid;
	wire [0 : 0]fork_43_out2_data;
	wire fork_43_out2_ready;
	wire fork_43_out2_valid;
	wire [0 : 0]fork_43_out3_data;
	wire fork_43_out3_ready;
	wire fork_43_out3_valid;

	wire cst_40_clk;
	wire cst_40_rst;
	wire [0 : 0]cst_40_in1_data;
	wire cst_40_in1_ready;
	wire cst_40_in1_valid;
	wire [0 : 0]cst_40_out1_data;
	wire cst_40_out1_ready;
	wire cst_40_out1_valid;

	wire phiC_30_clk;
	wire phiC_30_rst;
	wire [0 : 0]phiC_30_in1_data;
	wire phiC_30_in1_ready;
	wire phiC_30_in1_valid;
	wire [0 : 0]phiC_30_out1_data;
	wire phiC_30_out1_ready;
	wire phiC_30_out1_valid;

	wire forkC_65_clk;
	wire forkC_65_rst;
	wire [0 : 0]forkC_65_in1_data;
	wire forkC_65_in1_ready;
	wire forkC_65_in1_valid;
	wire [0 : 0]forkC_65_out1_data;
	wire forkC_65_out1_ready;
	wire forkC_65_out1_valid;
	wire [0 : 0]forkC_65_out2_data;
	wire forkC_65_out2_ready;
	wire forkC_65_out2_valid;

	wire branchC_52_clk;
	wire branchC_52_rst;
	wire [0 : 0]branchC_52_in1_data;
	wire branchC_52_in1_ready;
	wire branchC_52_in1_valid;
	wire [0 : 0]branchC_52_in2_data;
	wire branchC_52_in2_ready;
	wire branchC_52_in2_valid;
	wire [0 : 0]branchC_52_out1_data;
	wire branchC_52_out1_ready;
	wire branchC_52_out1_valid;
	wire [0 : 0]branchC_52_out2_data;
	wire branchC_52_out2_ready;
	wire branchC_52_out2_valid;

	wire source_15_clk;
	wire source_15_rst;
	wire [1 : 0]source_15_out1_data;
	wire source_15_out1_ready;
	wire source_15_out1_valid;

	wire source_16_clk;
	wire source_16_rst;
	wire [0 : 0]source_16_out1_data;
	wire source_16_out1_ready;
	wire source_16_out1_valid;

	wire source_17_clk;
	wire source_17_rst;
	wire [3 : 0]source_17_out1_data;
	wire source_17_out1_ready;
	wire source_17_out1_valid;

	wire phi_40_clk;
	wire phi_40_rst;
	wire [0 : 0]phi_40_in1_data;
	wire phi_40_in1_ready;
	wire phi_40_in1_valid;
	wire [3 : 0]phi_40_in2_data;
	wire phi_40_in2_ready;
	wire phi_40_in2_valid;
	wire [3 : 0]phi_40_in3_data;
	wire phi_40_in3_ready;
	wire phi_40_in3_valid;
	wire [3 : 0]phi_40_out1_data;
	wire phi_40_out1_ready;
	wire phi_40_out1_valid;

	wire cst_15_clk;
	wire cst_15_rst;
	wire [1 : 0]cst_15_in1_data;
	wire cst_15_in1_ready;
	wire cst_15_in1_valid;
	wire [1 : 0]cst_15_out1_data;
	wire cst_15_out1_ready;
	wire cst_15_out1_valid;

	wire shl_41_clk;
	wire shl_41_rst;
	wire [6 : 0]shl_41_in1_data;
	wire shl_41_in1_ready;
	wire shl_41_in1_valid;
	wire [6 : 0]shl_41_in2_data;
	wire shl_41_in2_ready;
	wire shl_41_in2_valid;
	wire [6 : 0]shl_41_out1_data;
	wire shl_41_out1_ready;
	wire shl_41_out1_valid;

	wire add_42_clk;
	wire add_42_rst;
	wire [7 : 0]add_42_in1_data;
	wire add_42_in1_ready;
	wire add_42_in1_valid;
	wire [7 : 0]add_42_in2_data;
	wire add_42_in2_ready;
	wire add_42_in2_valid;
	wire [7 : 0]add_42_out1_data;
	wire add_42_out1_ready;
	wire add_42_out1_valid;

	wire load_45_clk;
	wire load_45_rst;
	wire [31 : 0]load_45_in1_data;
	wire load_45_in1_ready;
	wire load_45_in1_valid;
	wire [7 : 0]load_45_in2_data;
	wire load_45_in2_ready;
	wire load_45_in2_valid;
	wire [31 : 0]load_45_out1_data;
	wire load_45_out1_ready;
	wire load_45_out1_valid;
	wire [7 : 0]load_45_out2_data;
	wire load_45_out2_ready;
	wire load_45_out2_valid;

	wire brCst_block9_clk;
	wire brCst_block9_rst;
	wire [0 : 0]brCst_block9_in1_data;
	wire brCst_block9_in1_ready;
	wire brCst_block9_in1_valid;
	wire [0 : 0]brCst_block9_out1_data;
	wire brCst_block9_out1_ready;
	wire brCst_block9_out1_valid;

	wire cst_16_clk;
	wire cst_16_rst;
	wire [0 : 0]cst_16_in1_data;
	wire cst_16_in1_ready;
	wire cst_16_in1_valid;
	wire [0 : 0]cst_16_out1_data;
	wire cst_16_out1_ready;
	wire cst_16_out1_valid;

	wire phi_n13_clk;
	wire phi_n13_rst;
	wire [3 : 0]phi_n13_in1_data;
	wire phi_n13_in1_ready;
	wire phi_n13_in1_valid;
	wire [3 : 0]phi_n13_in2_data;
	wire phi_n13_in2_ready;
	wire phi_n13_in2_valid;
	wire [3 : 0]phi_n13_out1_data;
	wire phi_n13_out1_ready;
	wire phi_n13_out1_valid;

	wire fork_6_clk;
	wire fork_6_rst;
	wire [3 : 0]fork_6_in1_data;
	wire fork_6_in1_ready;
	wire fork_6_in1_valid;
	wire [3 : 0]fork_6_out1_data;
	wire fork_6_out1_ready;
	wire fork_6_out1_valid;
	wire [3 : 0]fork_6_out2_data;
	wire fork_6_out2_ready;
	wire fork_6_out2_valid;

	wire fork_27_clk;
	wire fork_27_rst;
	wire [3 : 0]fork_27_in1_data;
	wire fork_27_in1_ready;
	wire fork_27_in1_valid;
	wire [3 : 0]fork_27_out1_data;
	wire fork_27_out1_ready;
	wire fork_27_out1_valid;
	wire [3 : 0]fork_27_out2_data;
	wire fork_27_out2_ready;
	wire fork_27_out2_valid;

	wire branch_17_clk;
	wire branch_17_rst;
	wire [31 : 0]branch_17_in1_data;
	wire branch_17_in1_ready;
	wire branch_17_in1_valid;
	wire [0 : 0]branch_17_in2_data;
	wire branch_17_in2_ready;
	wire branch_17_in2_valid;
	wire [31 : 0]branch_17_out1_data;
	wire branch_17_out1_ready;
	wire branch_17_out1_valid;
	wire [31 : 0]branch_17_out2_data;
	wire branch_17_out2_ready;
	wire branch_17_out2_valid;

	wire branch_18_clk;
	wire branch_18_rst;
	wire [0 : 0]branch_18_in1_data;
	wire branch_18_in1_ready;
	wire branch_18_in1_valid;
	wire [0 : 0]branch_18_in2_data;
	wire branch_18_in2_ready;
	wire branch_18_in2_valid;
	wire [0 : 0]branch_18_out1_data;
	wire branch_18_out1_ready;
	wire branch_18_out1_valid;
	wire [0 : 0]branch_18_out2_data;
	wire branch_18_out2_ready;
	wire branch_18_out2_valid;

	wire branch_19_clk;
	wire branch_19_rst;
	wire [3 : 0]branch_19_in1_data;
	wire branch_19_in1_ready;
	wire branch_19_in1_valid;
	wire [0 : 0]branch_19_in2_data;
	wire branch_19_in2_ready;
	wire branch_19_in2_valid;
	wire [3 : 0]branch_19_out1_data;
	wire branch_19_out1_ready;
	wire branch_19_out1_valid;
	wire [3 : 0]branch_19_out2_data;
	wire branch_19_out2_ready;
	wire branch_19_out2_valid;

	wire branch_20_clk;
	wire branch_20_rst;
	wire [3 : 0]branch_20_in1_data;
	wire branch_20_in1_ready;
	wire branch_20_in1_valid;
	wire [0 : 0]branch_20_in2_data;
	wire branch_20_in2_ready;
	wire branch_20_in2_valid;
	wire [3 : 0]branch_20_out1_data;
	wire branch_20_out1_ready;
	wire branch_20_out1_valid;
	wire [3 : 0]branch_20_out2_data;
	wire branch_20_out2_ready;
	wire branch_20_out2_valid;

	wire fork_41_clk;
	wire fork_41_rst;
	wire [0 : 0]fork_41_in1_data;
	wire fork_41_in1_ready;
	wire fork_41_in1_valid;
	wire [0 : 0]fork_41_out1_data;
	wire fork_41_out1_ready;
	wire fork_41_out1_valid;
	wire [0 : 0]fork_41_out2_data;
	wire fork_41_out2_ready;
	wire fork_41_out2_valid;
	wire [0 : 0]fork_41_out3_data;
	wire fork_41_out3_ready;
	wire fork_41_out3_valid;
	wire [0 : 0]fork_41_out4_data;
	wire fork_41_out4_ready;
	wire fork_41_out4_valid;
	wire [0 : 0]fork_41_out5_data;
	wire fork_41_out5_ready;
	wire fork_41_out5_valid;

	wire phiC_28_clk;
	wire phiC_28_rst;
	wire [0 : 0]phiC_28_in1_data;
	wire phiC_28_in1_ready;
	wire phiC_28_in1_valid;
	wire [0 : 0]phiC_28_in2_data;
	wire phiC_28_in2_ready;
	wire phiC_28_in2_valid;
	wire [0 : 0]phiC_28_out1_data;
	wire phiC_28_out1_ready;
	wire phiC_28_out1_valid;
	wire [0 : 0]phiC_28_out2_data;
	wire phiC_28_out2_ready;
	wire phiC_28_out2_valid;

	wire forkC_63_clk;
	wire forkC_63_rst;
	wire [0 : 0]forkC_63_in1_data;
	wire forkC_63_in1_ready;
	wire forkC_63_in1_valid;
	wire [0 : 0]forkC_63_out1_data;
	wire forkC_63_out1_ready;
	wire forkC_63_out1_valid;
	wire [0 : 0]forkC_63_out2_data;
	wire forkC_63_out2_ready;
	wire forkC_63_out2_valid;
	wire [0 : 0]forkC_63_out3_data;
	wire forkC_63_out3_ready;
	wire forkC_63_out3_valid;

	wire branchC_50_clk;
	wire branchC_50_rst;
	wire [0 : 0]branchC_50_in1_data;
	wire branchC_50_in1_ready;
	wire branchC_50_in1_valid;
	wire [0 : 0]branchC_50_in2_data;
	wire branchC_50_in2_ready;
	wire branchC_50_in2_valid;
	wire [0 : 0]branchC_50_out1_data;
	wire branchC_50_out1_ready;
	wire branchC_50_out1_valid;
	wire [0 : 0]branchC_50_out2_data;
	wire branchC_50_out2_ready;
	wire branchC_50_out2_valid;

	wire source_10_clk;
	wire source_10_rst;
	wire [1 : 0]source_10_out1_data;
	wire source_10_out1_ready;
	wire source_10_out1_valid;

	wire brCst_block7_clk;
	wire brCst_block7_rst;
	wire [0 : 0]brCst_block7_in1_data;
	wire brCst_block7_in1_ready;
	wire brCst_block7_in1_valid;
	wire [0 : 0]brCst_block7_out1_data;
	wire brCst_block7_out1_ready;
	wire brCst_block7_out1_valid;

	wire cst_13_clk;
	wire cst_13_rst;
	wire [0 : 0]cst_13_in1_data;
	wire cst_13_in1_ready;
	wire cst_13_in1_valid;
	wire [0 : 0]cst_13_out1_data;
	wire cst_13_out1_ready;
	wire cst_13_out1_valid;

	wire branch_14_clk;
	wire branch_14_rst;
	wire [0 : 0]branch_14_in1_data;
	wire branch_14_in1_ready;
	wire branch_14_in1_valid;
	wire [0 : 0]branch_14_in2_data;
	wire branch_14_in2_ready;
	wire branch_14_in2_valid;
	wire [0 : 0]branch_14_out1_data;
	wire branch_14_out1_ready;
	wire branch_14_out1_valid;
	wire [0 : 0]branch_14_out2_data;
	wire branch_14_out2_ready;
	wire branch_14_out2_valid;

	wire phiC_26_clk;
	wire phiC_26_rst;
	wire [0 : 0]phiC_26_in1_data;
	wire phiC_26_in1_ready;
	wire phiC_26_in1_valid;
	wire [0 : 0]phiC_26_out1_data;
	wire phiC_26_out1_ready;
	wire phiC_26_out1_valid;

	wire forkC_60_clk;
	wire forkC_60_rst;
	wire [0 : 0]forkC_60_in1_data;
	wire forkC_60_in1_ready;
	wire forkC_60_in1_valid;
	wire [0 : 0]forkC_60_out1_data;
	wire forkC_60_out1_ready;
	wire forkC_60_out1_valid;
	wire [0 : 0]forkC_60_out2_data;
	wire forkC_60_out2_ready;
	wire forkC_60_out2_valid;
	wire [0 : 0]forkC_60_out3_data;
	wire forkC_60_out3_ready;
	wire forkC_60_out3_valid;

	wire branchC_48_clk;
	wire branchC_48_rst;
	wire [0 : 0]branchC_48_in1_data;
	wire branchC_48_in1_ready;
	wire branchC_48_in1_valid;
	wire [0 : 0]branchC_48_in2_data;
	wire branchC_48_in2_ready;
	wire branchC_48_in2_valid;
	wire [0 : 0]branchC_48_out1_data;
	wire branchC_48_out1_ready;
	wire branchC_48_out1_valid;
	wire [0 : 0]branchC_48_out2_data;
	wire branchC_48_out2_ready;
	wire branchC_48_out2_valid;

	wire fork_61_clk;
	wire fork_61_rst;
	wire [0 : 0]fork_61_in1_data;
	wire fork_61_in1_ready;
	wire fork_61_in1_valid;
	wire [0 : 0]fork_61_out1_data;
	wire fork_61_out1_ready;
	wire fork_61_out1_valid;
	wire [0 : 0]fork_61_out2_data;
	wire fork_61_out2_ready;
	wire fork_61_out2_valid;

	wire brCst_block13_clk;
	wire brCst_block13_rst;
	wire [0 : 0]brCst_block13_in1_data;
	wire brCst_block13_in1_ready;
	wire brCst_block13_in1_valid;
	wire [0 : 0]brCst_block13_out1_data;
	wire brCst_block13_out1_ready;
	wire brCst_block13_out1_valid;

	wire cst_26_clk;
	wire cst_26_rst;
	wire [0 : 0]cst_26_in1_data;
	wire cst_26_in1_ready;
	wire cst_26_in1_valid;
	wire [0 : 0]cst_26_out1_data;
	wire cst_26_out1_ready;
	wire cst_26_out1_valid;

	wire branch_28_clk;
	wire branch_28_rst;
	wire [0 : 0]branch_28_in1_data;
	wire branch_28_in1_ready;
	wire branch_28_in1_valid;
	wire [0 : 0]branch_28_in2_data;
	wire branch_28_in2_ready;
	wire branch_28_in2_valid;
	wire [0 : 0]branch_28_out1_data;
	wire branch_28_out1_ready;
	wire branch_28_out1_valid;
	wire [0 : 0]branch_28_out2_data;
	wire branch_28_out2_ready;
	wire branch_28_out2_valid;

	wire phiC_32_clk;
	wire phiC_32_rst;
	wire [0 : 0]phiC_32_in1_data;
	wire phiC_32_in1_ready;
	wire phiC_32_in1_valid;
	wire [0 : 0]phiC_32_out1_data;
	wire phiC_32_out1_ready;
	wire phiC_32_out1_valid;

	wire forkC_68_clk;
	wire forkC_68_rst;
	wire [0 : 0]forkC_68_in1_data;
	wire forkC_68_in1_ready;
	wire forkC_68_in1_valid;
	wire [0 : 0]forkC_68_out1_data;
	wire forkC_68_out1_ready;
	wire forkC_68_out1_valid;
	wire [0 : 0]forkC_68_out2_data;
	wire forkC_68_out2_ready;
	wire forkC_68_out2_valid;
	wire [0 : 0]forkC_68_out3_data;
	wire forkC_68_out3_ready;
	wire forkC_68_out3_valid;

	wire branchC_54_clk;
	wire branchC_54_rst;
	wire [0 : 0]branchC_54_in1_data;
	wire branchC_54_in1_ready;
	wire branchC_54_in1_valid;
	wire [0 : 0]branchC_54_in2_data;
	wire branchC_54_in2_ready;
	wire branchC_54_in2_valid;
	wire [0 : 0]branchC_54_out1_data;
	wire branchC_54_out1_ready;
	wire branchC_54_out1_valid;
	wire [0 : 0]branchC_54_out2_data;
	wire branchC_54_out2_ready;
	wire branchC_54_out2_valid;

	wire fork_69_clk;
	wire fork_69_rst;
	wire [0 : 0]fork_69_in1_data;
	wire fork_69_in1_ready;
	wire fork_69_in1_valid;
	wire [0 : 0]fork_69_out1_data;
	wire fork_69_out1_ready;
	wire fork_69_out1_valid;
	wire [0 : 0]fork_69_out2_data;
	wire fork_69_out2_ready;
	wire fork_69_out2_valid;

	wire phi_75_clk;
	wire phi_75_rst;
	wire [0 : 0]phi_75_in1_data;
	wire phi_75_in1_ready;
	wire phi_75_in1_valid;
	wire [3 : 0]phi_75_in2_data;
	wire phi_75_in2_ready;
	wire phi_75_in2_valid;
	wire [3 : 0]phi_75_in3_data;
	wire phi_75_in3_ready;
	wire phi_75_in3_valid;
	wire [3 : 0]phi_75_out1_data;
	wire phi_75_out1_ready;
	wire phi_75_out1_valid;

	wire brCst_block14_clk;
	wire brCst_block14_rst;
	wire [0 : 0]brCst_block14_in1_data;
	wire brCst_block14_in1_ready;
	wire brCst_block14_in1_valid;
	wire [0 : 0]brCst_block14_out1_data;
	wire brCst_block14_out1_ready;
	wire brCst_block14_out1_valid;

	wire cst_27_clk;
	wire cst_27_rst;
	wire [0 : 0]cst_27_in1_data;
	wire cst_27_in1_ready;
	wire cst_27_in1_valid;
	wire [0 : 0]cst_27_out1_data;
	wire cst_27_out1_ready;
	wire cst_27_out1_valid;

	wire branch_29_clk;
	wire branch_29_rst;
	wire [0 : 0]branch_29_in1_data;
	wire branch_29_in1_ready;
	wire branch_29_in1_valid;
	wire [0 : 0]branch_29_in2_data;
	wire branch_29_in2_ready;
	wire branch_29_in2_valid;
	wire [0 : 0]branch_29_out1_data;
	wire branch_29_out1_ready;
	wire branch_29_out1_valid;
	wire [0 : 0]branch_29_out2_data;
	wire branch_29_out2_ready;
	wire branch_29_out2_valid;

	wire branch_30_clk;
	wire branch_30_rst;
	wire [3 : 0]branch_30_in1_data;
	wire branch_30_in1_ready;
	wire branch_30_in1_valid;
	wire [0 : 0]branch_30_in2_data;
	wire branch_30_in2_ready;
	wire branch_30_in2_valid;
	wire [3 : 0]branch_30_out1_data;
	wire branch_30_out1_ready;
	wire branch_30_out1_valid;
	wire [3 : 0]branch_30_out2_data;
	wire branch_30_out2_ready;
	wire branch_30_out2_valid;

	wire fork_46_clk;
	wire fork_46_rst;
	wire [0 : 0]fork_46_in1_data;
	wire fork_46_in1_ready;
	wire fork_46_in1_valid;
	wire [0 : 0]fork_46_out1_data;
	wire fork_46_out1_ready;
	wire fork_46_out1_valid;
	wire [0 : 0]fork_46_out2_data;
	wire fork_46_out2_ready;
	wire fork_46_out2_valid;
	wire [0 : 0]fork_46_out3_data;
	wire fork_46_out3_ready;
	wire fork_46_out3_valid;

	wire phiC_33_clk;
	wire phiC_33_rst;
	wire [0 : 0]phiC_33_in1_data;
	wire phiC_33_in1_ready;
	wire phiC_33_in1_valid;
	wire [0 : 0]phiC_33_in2_data;
	wire phiC_33_in2_ready;
	wire phiC_33_in2_valid;
	wire [0 : 0]phiC_33_out1_data;
	wire phiC_33_out1_ready;
	wire phiC_33_out1_valid;
	wire [0 : 0]phiC_33_out2_data;
	wire phiC_33_out2_ready;
	wire phiC_33_out2_valid;

	wire forkC_70_clk;
	wire forkC_70_rst;
	wire [0 : 0]forkC_70_in1_data;
	wire forkC_70_in1_ready;
	wire forkC_70_in1_valid;
	wire [0 : 0]forkC_70_out1_data;
	wire forkC_70_out1_ready;
	wire forkC_70_out1_valid;
	wire [0 : 0]forkC_70_out2_data;
	wire forkC_70_out2_ready;
	wire forkC_70_out2_valid;
	wire [0 : 0]forkC_70_out3_data;
	wire forkC_70_out3_ready;
	wire forkC_70_out3_valid;

	wire branchC_55_clk;
	wire branchC_55_rst;
	wire [0 : 0]branchC_55_in1_data;
	wire branchC_55_in1_ready;
	wire branchC_55_in1_valid;
	wire [0 : 0]branchC_55_in2_data;
	wire branchC_55_in2_ready;
	wire branchC_55_in2_valid;
	wire [0 : 0]branchC_55_out1_data;
	wire branchC_55_out1_ready;
	wire branchC_55_out1_valid;
	wire [0 : 0]branchC_55_out2_data;
	wire branchC_55_out2_ready;
	wire branchC_55_out2_valid;

	wire cst_37_clk;
	wire cst_37_rst;
	wire [0 : 0]cst_37_in1_data;
	wire cst_37_in1_ready;
	wire cst_37_in1_valid;
	wire [0 : 0]cst_37_out1_data;
	wire cst_37_out1_ready;
	wire cst_37_out1_valid;

	wire add_108_clk;
	wire add_108_rst;
	wire [3 : 0]add_108_in1_data;
	wire add_108_in1_ready;
	wire add_108_in1_valid;
	wire [3 : 0]add_108_in2_data;
	wire add_108_in2_ready;
	wire add_108_in2_valid;
	wire [3 : 0]add_108_out1_data;
	wire add_108_out1_ready;
	wire add_108_out1_valid;

	wire cst_38_clk;
	wire cst_38_rst;
	wire [3 : 0]cst_38_in1_data;
	wire cst_38_in1_ready;
	wire cst_38_in1_valid;
	wire [3 : 0]cst_38_out1_data;
	wire cst_38_out1_ready;
	wire cst_38_out1_valid;

	wire icmp_109_clk;
	wire icmp_109_rst;
	wire [3 : 0]icmp_109_in1_data;
	wire icmp_109_in1_ready;
	wire icmp_109_in1_valid;
	wire [3 : 0]icmp_109_in2_data;
	wire icmp_109_in2_ready;
	wire icmp_109_in2_valid;
	wire [0 : 0]icmp_109_out1_data;
	wire icmp_109_out1_ready;
	wire icmp_109_out1_valid;

	wire phi_n14_clk;
	wire phi_n14_rst;
	wire [3 : 0]phi_n14_in1_data;
	wire phi_n14_in1_ready;
	wire phi_n14_in1_valid;
	wire [3 : 0]phi_n14_out1_data;
	wire phi_n14_out1_ready;
	wire phi_n14_out1_valid;

	wire fork_17_clk;
	wire fork_17_rst;
	wire [3 : 0]fork_17_in1_data;
	wire fork_17_in1_ready;
	wire fork_17_in1_valid;
	wire [3 : 0]fork_17_out1_data;
	wire fork_17_out1_ready;
	wire fork_17_out1_valid;
	wire [3 : 0]fork_17_out2_data;
	wire fork_17_out2_ready;
	wire fork_17_out2_valid;

	wire branch_41_clk;
	wire branch_41_rst;
	wire [3 : 0]branch_41_in1_data;
	wire branch_41_in1_ready;
	wire branch_41_in1_valid;
	wire [0 : 0]branch_41_in2_data;
	wire branch_41_in2_ready;
	wire branch_41_in2_valid;
	wire [3 : 0]branch_41_out1_data;
	wire branch_41_out1_ready;
	wire branch_41_out1_valid;
	wire [3 : 0]branch_41_out2_data;
	wire branch_41_out2_ready;
	wire branch_41_out2_valid;

	wire phiC_37_clk;
	wire phiC_37_rst;
	wire [0 : 0]phiC_37_in1_data;
	wire phiC_37_in1_ready;
	wire phiC_37_in1_valid;
	wire [0 : 0]phiC_37_out1_data;
	wire phiC_37_out1_ready;
	wire phiC_37_out1_valid;

	wire branchC_59_clk;
	wire branchC_59_rst;
	wire [0 : 0]branchC_59_in1_data;
	wire branchC_59_in1_ready;
	wire branchC_59_in1_valid;
	wire [0 : 0]branchC_59_in2_data;
	wire branchC_59_in2_ready;
	wire branchC_59_in2_valid;
	wire [0 : 0]branchC_59_out1_data;
	wire branchC_59_out1_ready;
	wire branchC_59_out1_valid;
	wire [0 : 0]branchC_59_out2_data;
	wire branchC_59_out2_ready;
	wire branchC_59_out2_valid;

	wire fork_75_clk;
	wire fork_75_rst;
	wire [0 : 0]fork_75_in1_data;
	wire fork_75_in1_ready;
	wire fork_75_in1_valid;
	wire [0 : 0]fork_75_out1_data;
	wire fork_75_out1_ready;
	wire fork_75_out1_valid;
	wire [0 : 0]fork_75_out2_data;
	wire fork_75_out2_ready;
	wire fork_75_out2_valid;

	wire source_28_clk;
	wire source_28_rst;
	wire [0 : 0]source_28_out1_data;
	wire source_28_out1_ready;
	wire source_28_out1_valid;

	wire source_29_clk;
	wire source_29_rst;
	wire [3 : 0]source_29_out1_data;
	wire source_29_out1_ready;
	wire source_29_out1_valid;

	wire ret_0_clk;
	wire ret_0_rst;
	wire [0 : 0]ret_0_in1_data;
	wire ret_0_in1_ready;
	wire ret_0_in1_valid;
	wire [0 : 0]ret_0_out1_data;
	wire ret_0_out1_ready;
	wire ret_0_out1_valid;

	wire end_0_clk;
	wire end_0_rst;
	wire [0 : 0]end_0_in1_data;
	wire end_0_in1_ready;
	wire end_0_in1_valid;
	wire [0 : 0]end_0_in2_data;
	wire end_0_in2_ready;
	wire end_0_in2_valid;
	wire [0 : 0]end_0_in3_data;
	wire end_0_in3_ready;
	wire end_0_in3_valid;
	wire [0 : 0]end_0_in4_data;
	wire end_0_in4_ready;
	wire end_0_in4_valid;
	wire [0 : 0]end_0_in5_data;
	wire end_0_in5_ready;
	wire end_0_in5_valid;
	wire [0 : 0]end_0_in6_data;
	wire end_0_in6_ready;
	wire end_0_in6_valid;
	wire [0 : 0]end_0_in7_data;
	wire end_0_in7_ready;
	wire end_0_in7_valid;
	wire [0 : 0]end_0_in8_data;
	wire end_0_in8_ready;
	wire end_0_in8_valid;
	wire [0 : 0]end_0_out1_data;
	wire end_0_out1_ready;
	wire end_0_out1_valid;

	wire phiC_38_clk;
	wire phiC_38_rst;
	wire [0 : 0]phiC_38_in1_data;
	wire phiC_38_in1_ready;
	wire phiC_38_in1_valid;
	wire [0 : 0]phiC_38_out1_data;
	wire phiC_38_out1_ready;
	wire phiC_38_out1_valid;

	wire cst_24_clk;
	wire cst_24_rst;
	wire [0 : 0]cst_24_in1_data;
	wire cst_24_in1_ready;
	wire cst_24_in1_valid;
	wire [0 : 0]cst_24_out1_data;
	wire cst_24_out1_ready;
	wire cst_24_out1_valid;

	wire add_71_clk;
	wire add_71_rst;
	wire [3 : 0]add_71_in1_data;
	wire add_71_in1_ready;
	wire add_71_in1_valid;
	wire [3 : 0]add_71_in2_data;
	wire add_71_in2_ready;
	wire add_71_in2_valid;
	wire [3 : 0]add_71_out1_data;
	wire add_71_out1_ready;
	wire add_71_out1_valid;

	wire cst_25_clk;
	wire cst_25_rst;
	wire [3 : 0]cst_25_in1_data;
	wire cst_25_in1_ready;
	wire cst_25_in1_valid;
	wire [3 : 0]cst_25_out1_data;
	wire cst_25_out1_ready;
	wire cst_25_out1_valid;

	wire icmp_72_clk;
	wire icmp_72_rst;
	wire [3 : 0]icmp_72_in1_data;
	wire icmp_72_in1_ready;
	wire icmp_72_in1_valid;
	wire [3 : 0]icmp_72_in2_data;
	wire icmp_72_in2_ready;
	wire icmp_72_in2_valid;
	wire [0 : 0]icmp_72_out1_data;
	wire icmp_72_out1_ready;
	wire icmp_72_out1_valid;

	wire phi_n12_clk;
	wire phi_n12_rst;
	wire [3 : 0]phi_n12_in1_data;
	wire phi_n12_in1_ready;
	wire phi_n12_in1_valid;
	wire [3 : 0]phi_n12_out1_data;
	wire phi_n12_out1_ready;
	wire phi_n12_out1_valid;

	wire fork_11_clk;
	wire fork_11_rst;
	wire [3 : 0]fork_11_in1_data;
	wire fork_11_in1_ready;
	wire fork_11_in1_valid;
	wire [3 : 0]fork_11_out1_data;
	wire fork_11_out1_ready;
	wire fork_11_out1_valid;
	wire [3 : 0]fork_11_out2_data;
	wire fork_11_out2_ready;
	wire fork_11_out2_valid;

	wire branch_27_clk;
	wire branch_27_rst;
	wire [3 : 0]branch_27_in1_data;
	wire branch_27_in1_ready;
	wire branch_27_in1_valid;
	wire [0 : 0]branch_27_in2_data;
	wire branch_27_in2_ready;
	wire branch_27_in2_valid;
	wire [3 : 0]branch_27_out1_data;
	wire branch_27_out1_ready;
	wire branch_27_out1_valid;
	wire [3 : 0]branch_27_out2_data;
	wire branch_27_out2_ready;
	wire branch_27_out2_valid;

	wire phiC_31_clk;
	wire phiC_31_rst;
	wire [0 : 0]phiC_31_in1_data;
	wire phiC_31_in1_ready;
	wire phiC_31_in1_valid;
	wire [0 : 0]phiC_31_out1_data;
	wire phiC_31_out1_ready;
	wire phiC_31_out1_valid;

	wire branchC_53_clk;
	wire branchC_53_rst;
	wire [0 : 0]branchC_53_in1_data;
	wire branchC_53_in1_ready;
	wire branchC_53_in1_valid;
	wire [0 : 0]branchC_53_in2_data;
	wire branchC_53_in2_ready;
	wire branchC_53_in2_valid;
	wire [0 : 0]branchC_53_out1_data;
	wire branchC_53_out1_ready;
	wire branchC_53_out1_valid;
	wire [0 : 0]branchC_53_out2_data;
	wire branchC_53_out2_ready;
	wire branchC_53_out2_valid;

	wire fork_67_clk;
	wire fork_67_rst;
	wire [0 : 0]fork_67_in1_data;
	wire fork_67_in1_ready;
	wire fork_67_in1_valid;
	wire [0 : 0]fork_67_out1_data;
	wire fork_67_out1_ready;
	wire fork_67_out1_valid;
	wire [0 : 0]fork_67_out2_data;
	wire fork_67_out2_ready;
	wire fork_67_out2_valid;

	wire source_18_clk;
	wire source_18_rst;
	wire [0 : 0]source_18_out1_data;
	wire source_18_out1_ready;
	wire source_18_out1_valid;

	wire source_19_clk;
	wire source_19_rst;
	wire [3 : 0]source_19_out1_data;
	wire source_19_out1_ready;
	wire source_19_out1_valid;

	wire phi_47_clk;
	wire phi_47_rst;
	wire [0 : 0]phi_47_in1_data;
	wire phi_47_in1_ready;
	wire phi_47_in1_valid;
	wire [31 : 0]phi_47_in2_data;
	wire phi_47_in2_ready;
	wire phi_47_in2_valid;
	wire [31 : 0]phi_47_in3_data;
	wire phi_47_in3_ready;
	wire phi_47_in3_valid;
	wire [31 : 0]phi_47_out1_data;
	wire phi_47_out1_ready;
	wire phi_47_out1_valid;

	wire phi_48_clk;
	wire phi_48_rst;
	wire [0 : 0]phi_48_in1_data;
	wire phi_48_in1_ready;
	wire phi_48_in1_valid;
	wire [3 : 0]phi_48_in2_data;
	wire phi_48_in2_ready;
	wire phi_48_in2_valid;
	wire [3 : 0]phi_48_in3_data;
	wire phi_48_in3_ready;
	wire phi_48_in3_valid;
	wire [3 : 0]phi_48_out1_data;
	wire phi_48_out1_ready;
	wire phi_48_out1_valid;

	wire cst_17_clk;
	wire cst_17_rst;
	wire [1 : 0]cst_17_in1_data;
	wire cst_17_in1_ready;
	wire cst_17_in1_valid;
	wire [1 : 0]cst_17_out1_data;
	wire cst_17_out1_ready;
	wire cst_17_out1_valid;

	wire shl_49_clk;
	wire shl_49_rst;
	wire [6 : 0]shl_49_in1_data;
	wire shl_49_in1_ready;
	wire shl_49_in1_valid;
	wire [6 : 0]shl_49_in2_data;
	wire shl_49_in2_ready;
	wire shl_49_in2_valid;
	wire [6 : 0]shl_49_out1_data;
	wire shl_49_out1_ready;
	wire shl_49_out1_valid;

	wire add_50_clk;
	wire add_50_rst;
	wire [7 : 0]add_50_in1_data;
	wire add_50_in1_ready;
	wire add_50_in1_valid;
	wire [7 : 0]add_50_in2_data;
	wire add_50_in2_ready;
	wire add_50_in2_valid;
	wire [7 : 0]add_50_out1_data;
	wire add_50_out1_ready;
	wire add_50_out1_valid;

	wire load_53_clk;
	wire load_53_rst;
	wire [31 : 0]load_53_in1_data;
	wire load_53_in1_ready;
	wire load_53_in1_valid;
	wire [7 : 0]load_53_in2_data;
	wire load_53_in2_ready;
	wire load_53_in2_valid;
	wire [31 : 0]load_53_out1_data;
	wire load_53_out1_ready;
	wire load_53_out1_valid;
	wire [7 : 0]load_53_out2_data;
	wire load_53_out2_ready;
	wire load_53_out2_valid;

	wire cst_18_clk;
	wire cst_18_rst;
	wire [1 : 0]cst_18_in1_data;
	wire cst_18_in1_ready;
	wire cst_18_in1_valid;
	wire [1 : 0]cst_18_out1_data;
	wire cst_18_out1_ready;
	wire cst_18_out1_valid;

	wire shl_54_clk;
	wire shl_54_rst;
	wire [6 : 0]shl_54_in1_data;
	wire shl_54_in1_ready;
	wire shl_54_in1_valid;
	wire [6 : 0]shl_54_in2_data;
	wire shl_54_in2_ready;
	wire shl_54_in2_valid;
	wire [6 : 0]shl_54_out1_data;
	wire shl_54_out1_ready;
	wire shl_54_out1_valid;

	wire add_55_clk;
	wire add_55_rst;
	wire [7 : 0]add_55_in1_data;
	wire add_55_in1_ready;
	wire add_55_in1_valid;
	wire [7 : 0]add_55_in2_data;
	wire add_55_in2_ready;
	wire add_55_in2_valid;
	wire [7 : 0]add_55_out1_data;
	wire add_55_out1_ready;
	wire add_55_out1_valid;

	wire load_58_clk;
	wire load_58_rst;
	wire [31 : 0]load_58_in1_data;
	wire load_58_in1_ready;
	wire load_58_in1_valid;
	wire [7 : 0]load_58_in2_data;
	wire load_58_in2_ready;
	wire load_58_in2_valid;
	wire [31 : 0]load_58_out1_data;
	wire load_58_out1_ready;
	wire load_58_out1_valid;
	wire [7 : 0]load_58_out2_data;
	wire load_58_out2_ready;
	wire load_58_out2_valid;

	wire cst_19_clk;
	wire cst_19_rst;
	wire [0 : 0]cst_19_in1_data;
	wire cst_19_in1_ready;
	wire cst_19_in1_valid;
	wire [0 : 0]cst_19_out1_data;
	wire cst_19_out1_ready;
	wire cst_19_out1_valid;

	wire add_61_clk;
	wire add_61_rst;
	wire [3 : 0]add_61_in1_data;
	wire add_61_in1_ready;
	wire add_61_in1_valid;
	wire [3 : 0]add_61_in2_data;
	wire add_61_in2_ready;
	wire add_61_in2_valid;
	wire [3 : 0]add_61_out1_data;
	wire add_61_out1_ready;
	wire add_61_out1_valid;

	wire cst_20_clk;
	wire cst_20_rst;
	wire [3 : 0]cst_20_in1_data;
	wire cst_20_in1_ready;
	wire cst_20_in1_valid;
	wire [3 : 0]cst_20_out1_data;
	wire cst_20_out1_ready;
	wire cst_20_out1_valid;

	wire icmp_62_clk;
	wire icmp_62_rst;
	wire [3 : 0]icmp_62_in1_data;
	wire icmp_62_in1_ready;
	wire icmp_62_in1_valid;
	wire [3 : 0]icmp_62_in2_data;
	wire icmp_62_in2_ready;
	wire icmp_62_in2_valid;
	wire [0 : 0]icmp_62_out1_data;
	wire icmp_62_out1_ready;
	wire icmp_62_out1_valid;

	wire phi_n10_clk;
	wire phi_n10_rst;
	wire [3 : 0]phi_n10_in1_data;
	wire phi_n10_in1_ready;
	wire phi_n10_in1_valid;
	wire [3 : 0]phi_n10_in2_data;
	wire phi_n10_in2_ready;
	wire phi_n10_in2_valid;
	wire [3 : 0]phi_n10_out1_data;
	wire phi_n10_out1_ready;
	wire phi_n10_out1_valid;

	wire phi_n11_clk;
	wire phi_n11_rst;
	wire [3 : 0]phi_n11_in1_data;
	wire phi_n11_in1_ready;
	wire phi_n11_in1_valid;
	wire [3 : 0]phi_n11_in2_data;
	wire phi_n11_in2_ready;
	wire phi_n11_in2_valid;
	wire [3 : 0]phi_n11_out1_data;
	wire phi_n11_out1_ready;
	wire phi_n11_out1_valid;

	wire fork_7_clk;
	wire fork_7_rst;
	wire [3 : 0]fork_7_in1_data;
	wire fork_7_in1_ready;
	wire fork_7_in1_valid;
	wire [3 : 0]fork_7_out1_data;
	wire fork_7_out1_ready;
	wire fork_7_out1_valid;
	wire [3 : 0]fork_7_out2_data;
	wire fork_7_out2_ready;
	wire fork_7_out2_valid;
	wire [3 : 0]fork_7_out3_data;
	wire fork_7_out3_ready;
	wire fork_7_out3_valid;

	wire fork_9_clk;
	wire fork_9_rst;
	wire [3 : 0]fork_9_in1_data;
	wire fork_9_in1_ready;
	wire fork_9_in1_valid;
	wire [3 : 0]fork_9_out1_data;
	wire fork_9_out1_ready;
	wire fork_9_out1_valid;
	wire [3 : 0]fork_9_out2_data;
	wire fork_9_out2_ready;
	wire fork_9_out2_valid;

	wire fork_25_clk;
	wire fork_25_rst;
	wire [3 : 0]fork_25_in1_data;
	wire fork_25_in1_ready;
	wire fork_25_in1_valid;
	wire [3 : 0]fork_25_out1_data;
	wire fork_25_out1_ready;
	wire fork_25_out1_valid;
	wire [3 : 0]fork_25_out2_data;
	wire fork_25_out2_ready;
	wire fork_25_out2_valid;

	wire fork_26_clk;
	wire fork_26_rst;
	wire [3 : 0]fork_26_in1_data;
	wire fork_26_in1_ready;
	wire fork_26_in1_valid;
	wire [3 : 0]fork_26_out1_data;
	wire fork_26_out1_ready;
	wire fork_26_out1_valid;
	wire [3 : 0]fork_26_out2_data;
	wire fork_26_out2_ready;
	wire fork_26_out2_valid;

	wire branch_21_clk;
	wire branch_21_rst;
	wire [31 : 0]branch_21_in1_data;
	wire branch_21_in1_ready;
	wire branch_21_in1_valid;
	wire [0 : 0]branch_21_in2_data;
	wire branch_21_in2_ready;
	wire branch_21_in2_valid;
	wire [31 : 0]branch_21_out1_data;
	wire branch_21_out1_ready;
	wire branch_21_out1_valid;
	wire [31 : 0]branch_21_out2_data;
	wire branch_21_out2_ready;
	wire branch_21_out2_valid;

	wire branch_22_clk;
	wire branch_22_rst;
	wire [3 : 0]branch_22_in1_data;
	wire branch_22_in1_ready;
	wire branch_22_in1_valid;
	wire [0 : 0]branch_22_in2_data;
	wire branch_22_in2_ready;
	wire branch_22_in2_valid;
	wire [3 : 0]branch_22_out1_data;
	wire branch_22_out1_ready;
	wire branch_22_out1_valid;
	wire [3 : 0]branch_22_out2_data;
	wire branch_22_out2_ready;
	wire branch_22_out2_valid;

	wire branch_23_clk;
	wire branch_23_rst;
	wire [3 : 0]branch_23_in1_data;
	wire branch_23_in1_ready;
	wire branch_23_in1_valid;
	wire [0 : 0]branch_23_in2_data;
	wire branch_23_in2_ready;
	wire branch_23_in2_valid;
	wire [3 : 0]branch_23_out1_data;
	wire branch_23_out1_ready;
	wire branch_23_out1_valid;
	wire [3 : 0]branch_23_out2_data;
	wire branch_23_out2_ready;
	wire branch_23_out2_valid;

	wire branch_24_clk;
	wire branch_24_rst;
	wire [3 : 0]branch_24_in1_data;
	wire branch_24_in1_ready;
	wire branch_24_in1_valid;
	wire [0 : 0]branch_24_in2_data;
	wire branch_24_in2_ready;
	wire branch_24_in2_valid;
	wire [3 : 0]branch_24_out1_data;
	wire branch_24_out1_ready;
	wire branch_24_out1_valid;
	wire [3 : 0]branch_24_out2_data;
	wire branch_24_out2_ready;
	wire branch_24_out2_valid;

	wire fork_42_clk;
	wire fork_42_rst;
	wire [0 : 0]fork_42_in1_data;
	wire fork_42_in1_ready;
	wire fork_42_in1_valid;
	wire [0 : 0]fork_42_out1_data;
	wire fork_42_out1_ready;
	wire fork_42_out1_valid;
	wire [0 : 0]fork_42_out2_data;
	wire fork_42_out2_ready;
	wire fork_42_out2_valid;
	wire [0 : 0]fork_42_out3_data;
	wire fork_42_out3_ready;
	wire fork_42_out3_valid;
	wire [0 : 0]fork_42_out4_data;
	wire fork_42_out4_ready;
	wire fork_42_out4_valid;
	wire [0 : 0]fork_42_out5_data;
	wire fork_42_out5_ready;
	wire fork_42_out5_valid;

	wire phiC_29_clk;
	wire phiC_29_rst;
	wire [0 : 0]phiC_29_in1_data;
	wire phiC_29_in1_ready;
	wire phiC_29_in1_valid;
	wire [0 : 0]phiC_29_in2_data;
	wire phiC_29_in2_ready;
	wire phiC_29_in2_valid;
	wire [0 : 0]phiC_29_out1_data;
	wire phiC_29_out1_ready;
	wire phiC_29_out1_valid;
	wire [0 : 0]phiC_29_out2_data;
	wire phiC_29_out2_ready;
	wire phiC_29_out2_valid;

	wire branchC_51_clk;
	wire branchC_51_rst;
	wire [0 : 0]branchC_51_in1_data;
	wire branchC_51_in1_ready;
	wire branchC_51_in1_valid;
	wire [0 : 0]branchC_51_in2_data;
	wire branchC_51_in2_ready;
	wire branchC_51_in2_valid;
	wire [0 : 0]branchC_51_out1_data;
	wire branchC_51_out1_ready;
	wire branchC_51_out1_valid;
	wire [0 : 0]branchC_51_out2_data;
	wire branchC_51_out2_ready;
	wire branchC_51_out2_valid;

	wire source_11_clk;
	wire source_11_rst;
	wire [1 : 0]source_11_out1_data;
	wire source_11_out1_ready;
	wire source_11_out1_valid;

	wire source_12_clk;
	wire source_12_rst;
	wire [1 : 0]source_12_out1_data;
	wire source_12_out1_ready;
	wire source_12_out1_valid;

	wire source_13_clk;
	wire source_13_rst;
	wire [0 : 0]source_13_out1_data;
	wire source_13_out1_ready;
	wire source_13_out1_valid;

	wire source_14_clk;
	wire source_14_rst;
	wire [3 : 0]source_14_out1_data;
	wire source_14_out1_ready;
	wire source_14_out1_valid;

	wire fork_82_clk;
	wire fork_82_rst;
	wire [0 : 0]fork_82_in1_data;
	wire fork_82_in1_ready;
	wire fork_82_in1_valid;
	wire [0 : 0]fork_82_out1_data;
	wire fork_82_out1_ready;
	wire fork_82_out1_valid;
	wire [0 : 0]fork_82_out2_data;
	wire fork_82_out2_ready;
	wire fork_82_out2_valid;

	wire phi_10_clk;
	wire phi_10_rst;
	wire [0 : 0]phi_10_in1_data;
	wire phi_10_in1_ready;
	wire phi_10_in1_valid;
	wire [31 : 0]phi_10_in2_data;
	wire phi_10_in2_ready;
	wire phi_10_in2_valid;
	wire [31 : 0]phi_10_in3_data;
	wire phi_10_in3_ready;
	wire phi_10_in3_valid;
	wire [31 : 0]phi_10_out1_data;
	wire phi_10_out1_ready;
	wire phi_10_out1_valid;

	wire phi_11_clk;
	wire phi_11_rst;
	wire [0 : 0]phi_11_in1_data;
	wire phi_11_in1_ready;
	wire phi_11_in1_valid;
	wire [3 : 0]phi_11_in2_data;
	wire phi_11_in2_ready;
	wire phi_11_in2_valid;
	wire [3 : 0]phi_11_in3_data;
	wire phi_11_in3_ready;
	wire phi_11_in3_valid;
	wire [3 : 0]phi_11_out1_data;
	wire phi_11_out1_ready;
	wire phi_11_out1_valid;

	wire cst_4_clk;
	wire cst_4_rst;
	wire [1 : 0]cst_4_in1_data;
	wire cst_4_in1_ready;
	wire cst_4_in1_valid;
	wire [1 : 0]cst_4_out1_data;
	wire cst_4_out1_ready;
	wire cst_4_out1_valid;

	wire shl_12_clk;
	wire shl_12_rst;
	wire [6 : 0]shl_12_in1_data;
	wire shl_12_in1_ready;
	wire shl_12_in1_valid;
	wire [6 : 0]shl_12_in2_data;
	wire shl_12_in2_ready;
	wire shl_12_in2_valid;
	wire [6 : 0]shl_12_out1_data;
	wire shl_12_out1_ready;
	wire shl_12_out1_valid;

	wire add_13_clk;
	wire add_13_rst;
	wire [7 : 0]add_13_in1_data;
	wire add_13_in1_ready;
	wire add_13_in1_valid;
	wire [7 : 0]add_13_in2_data;
	wire add_13_in2_ready;
	wire add_13_in2_valid;
	wire [7 : 0]add_13_out1_data;
	wire add_13_out1_ready;
	wire add_13_out1_valid;

	wire load_16_clk;
	wire load_16_rst;
	wire [31 : 0]load_16_in1_data;
	wire load_16_in1_ready;
	wire load_16_in1_valid;
	wire [7 : 0]load_16_in2_data;
	wire load_16_in2_ready;
	wire load_16_in2_valid;
	wire [31 : 0]load_16_out1_data;
	wire load_16_out1_ready;
	wire load_16_out1_valid;
	wire [7 : 0]load_16_out2_data;
	wire load_16_out2_ready;
	wire load_16_out2_valid;

	wire cst_5_clk;
	wire cst_5_rst;
	wire [1 : 0]cst_5_in1_data;
	wire cst_5_in1_ready;
	wire cst_5_in1_valid;
	wire [1 : 0]cst_5_out1_data;
	wire cst_5_out1_ready;
	wire cst_5_out1_valid;

	wire shl_17_clk;
	wire shl_17_rst;
	wire [6 : 0]shl_17_in1_data;
	wire shl_17_in1_ready;
	wire shl_17_in1_valid;
	wire [6 : 0]shl_17_in2_data;
	wire shl_17_in2_ready;
	wire shl_17_in2_valid;
	wire [6 : 0]shl_17_out1_data;
	wire shl_17_out1_ready;
	wire shl_17_out1_valid;

	wire add_18_clk;
	wire add_18_rst;
	wire [7 : 0]add_18_in1_data;
	wire add_18_in1_ready;
	wire add_18_in1_valid;
	wire [7 : 0]add_18_in2_data;
	wire add_18_in2_ready;
	wire add_18_in2_valid;
	wire [7 : 0]add_18_out1_data;
	wire add_18_out1_ready;
	wire add_18_out1_valid;

	wire load_21_clk;
	wire load_21_rst;
	wire [31 : 0]load_21_in1_data;
	wire load_21_in1_ready;
	wire load_21_in1_valid;
	wire [7 : 0]load_21_in2_data;
	wire load_21_in2_ready;
	wire load_21_in2_valid;
	wire [31 : 0]load_21_out1_data;
	wire load_21_out1_ready;
	wire load_21_out1_valid;
	wire [7 : 0]load_21_out2_data;
	wire load_21_out2_ready;
	wire load_21_out2_valid;

	wire cst_6_clk;
	wire cst_6_rst;
	wire [0 : 0]cst_6_in1_data;
	wire cst_6_in1_ready;
	wire cst_6_in1_valid;
	wire [0 : 0]cst_6_out1_data;
	wire cst_6_out1_ready;
	wire cst_6_out1_valid;

	wire add_24_clk;
	wire add_24_rst;
	wire [3 : 0]add_24_in1_data;
	wire add_24_in1_ready;
	wire add_24_in1_valid;
	wire [3 : 0]add_24_in2_data;
	wire add_24_in2_ready;
	wire add_24_in2_valid;
	wire [3 : 0]add_24_out1_data;
	wire add_24_out1_ready;
	wire add_24_out1_valid;

	wire cst_7_clk;
	wire cst_7_rst;
	wire [3 : 0]cst_7_in1_data;
	wire cst_7_in1_ready;
	wire cst_7_in1_valid;
	wire [3 : 0]cst_7_out1_data;
	wire cst_7_out1_ready;
	wire cst_7_out1_valid;

	wire icmp_25_clk;
	wire icmp_25_rst;
	wire [3 : 0]icmp_25_in1_data;
	wire icmp_25_in1_ready;
	wire icmp_25_in1_valid;
	wire [3 : 0]icmp_25_in2_data;
	wire icmp_25_in2_ready;
	wire icmp_25_in2_valid;
	wire [0 : 0]icmp_25_out1_data;
	wire icmp_25_out1_ready;
	wire icmp_25_out1_valid;

	wire phi_n8_clk;
	wire phi_n8_rst;
	wire [3 : 0]phi_n8_in1_data;
	wire phi_n8_in1_ready;
	wire phi_n8_in1_valid;
	wire [3 : 0]phi_n8_in2_data;
	wire phi_n8_in2_ready;
	wire phi_n8_in2_valid;
	wire [3 : 0]phi_n8_out1_data;
	wire phi_n8_out1_ready;
	wire phi_n8_out1_valid;

	wire phi_n9_clk;
	wire phi_n9_rst;
	wire [3 : 0]phi_n9_in1_data;
	wire phi_n9_in1_ready;
	wire phi_n9_in1_valid;
	wire [3 : 0]phi_n9_in2_data;
	wire phi_n9_in2_ready;
	wire phi_n9_in2_valid;
	wire [3 : 0]phi_n9_out1_data;
	wire phi_n9_out1_ready;
	wire phi_n9_out1_valid;

	wire fork_1_clk;
	wire fork_1_rst;
	wire [3 : 0]fork_1_in1_data;
	wire fork_1_in1_ready;
	wire fork_1_in1_valid;
	wire [3 : 0]fork_1_out1_data;
	wire fork_1_out1_ready;
	wire fork_1_out1_valid;
	wire [3 : 0]fork_1_out2_data;
	wire fork_1_out2_ready;
	wire fork_1_out2_valid;
	wire [3 : 0]fork_1_out3_data;
	wire fork_1_out3_ready;
	wire fork_1_out3_valid;

	wire fork_3_clk;
	wire fork_3_rst;
	wire [3 : 0]fork_3_in1_data;
	wire fork_3_in1_ready;
	wire fork_3_in1_valid;
	wire [3 : 0]fork_3_out1_data;
	wire fork_3_out1_ready;
	wire fork_3_out1_valid;
	wire [3 : 0]fork_3_out2_data;
	wire fork_3_out2_ready;
	wire fork_3_out2_valid;

	wire fork_23_clk;
	wire fork_23_rst;
	wire [3 : 0]fork_23_in1_data;
	wire fork_23_in1_ready;
	wire fork_23_in1_valid;
	wire [3 : 0]fork_23_out1_data;
	wire fork_23_out1_ready;
	wire fork_23_out1_valid;
	wire [3 : 0]fork_23_out2_data;
	wire fork_23_out2_ready;
	wire fork_23_out2_valid;

	wire fork_24_clk;
	wire fork_24_rst;
	wire [3 : 0]fork_24_in1_data;
	wire fork_24_in1_ready;
	wire fork_24_in1_valid;
	wire [3 : 0]fork_24_out1_data;
	wire fork_24_out1_ready;
	wire fork_24_out1_valid;
	wire [3 : 0]fork_24_out2_data;
	wire fork_24_out2_ready;
	wire fork_24_out2_valid;

	wire branch_7_clk;
	wire branch_7_rst;
	wire [31 : 0]branch_7_in1_data;
	wire branch_7_in1_ready;
	wire branch_7_in1_valid;
	wire [0 : 0]branch_7_in2_data;
	wire branch_7_in2_ready;
	wire branch_7_in2_valid;
	wire [31 : 0]branch_7_out1_data;
	wire branch_7_out1_ready;
	wire branch_7_out1_valid;
	wire [31 : 0]branch_7_out2_data;
	wire branch_7_out2_ready;
	wire branch_7_out2_valid;

	wire branch_8_clk;
	wire branch_8_rst;
	wire [3 : 0]branch_8_in1_data;
	wire branch_8_in1_ready;
	wire branch_8_in1_valid;
	wire [0 : 0]branch_8_in2_data;
	wire branch_8_in2_ready;
	wire branch_8_in2_valid;
	wire [3 : 0]branch_8_out1_data;
	wire branch_8_out1_ready;
	wire branch_8_out1_valid;
	wire [3 : 0]branch_8_out2_data;
	wire branch_8_out2_ready;
	wire branch_8_out2_valid;

	wire branch_9_clk;
	wire branch_9_rst;
	wire [3 : 0]branch_9_in1_data;
	wire branch_9_in1_ready;
	wire branch_9_in1_valid;
	wire [0 : 0]branch_9_in2_data;
	wire branch_9_in2_ready;
	wire branch_9_in2_valid;
	wire [3 : 0]branch_9_out1_data;
	wire branch_9_out1_ready;
	wire branch_9_out1_valid;
	wire [3 : 0]branch_9_out2_data;
	wire branch_9_out2_ready;
	wire branch_9_out2_valid;

	wire branch_10_clk;
	wire branch_10_rst;
	wire [3 : 0]branch_10_in1_data;
	wire branch_10_in1_ready;
	wire branch_10_in1_valid;
	wire [0 : 0]branch_10_in2_data;
	wire branch_10_in2_ready;
	wire branch_10_in2_valid;
	wire [3 : 0]branch_10_out1_data;
	wire branch_10_out1_ready;
	wire branch_10_out1_valid;
	wire [3 : 0]branch_10_out2_data;
	wire branch_10_out2_ready;
	wire branch_10_out2_valid;

	wire fork_36_clk;
	wire fork_36_rst;
	wire [0 : 0]fork_36_in1_data;
	wire fork_36_in1_ready;
	wire fork_36_in1_valid;
	wire [0 : 0]fork_36_out1_data;
	wire fork_36_out1_ready;
	wire fork_36_out1_valid;
	wire [0 : 0]fork_36_out2_data;
	wire fork_36_out2_ready;
	wire fork_36_out2_valid;
	wire [0 : 0]fork_36_out3_data;
	wire fork_36_out3_ready;
	wire fork_36_out3_valid;
	wire [0 : 0]fork_36_out4_data;
	wire fork_36_out4_ready;
	wire fork_36_out4_valid;
	wire [0 : 0]fork_36_out5_data;
	wire fork_36_out5_ready;
	wire fork_36_out5_valid;

	wire phiC_23_clk;
	wire phiC_23_rst;
	wire [0 : 0]phiC_23_in1_data;
	wire phiC_23_in1_ready;
	wire phiC_23_in1_valid;
	wire [0 : 0]phiC_23_in2_data;
	wire phiC_23_in2_ready;
	wire phiC_23_in2_valid;
	wire [0 : 0]phiC_23_out1_data;
	wire phiC_23_out1_ready;
	wire phiC_23_out1_valid;
	wire [0 : 0]phiC_23_out2_data;
	wire phiC_23_out2_ready;
	wire phiC_23_out2_valid;

	wire branchC_45_clk;
	wire branchC_45_rst;
	wire [0 : 0]branchC_45_in1_data;
	wire branchC_45_in1_ready;
	wire branchC_45_in1_valid;
	wire [0 : 0]branchC_45_in2_data;
	wire branchC_45_in2_ready;
	wire branchC_45_in2_valid;
	wire [0 : 0]branchC_45_out1_data;
	wire branchC_45_out1_ready;
	wire branchC_45_out1_valid;
	wire [0 : 0]branchC_45_out2_data;
	wire branchC_45_out2_ready;
	wire branchC_45_out2_valid;

	wire source_1_clk;
	wire source_1_rst;
	wire [1 : 0]source_1_out1_data;
	wire source_1_out1_ready;
	wire source_1_out1_valid;

	wire source_2_clk;
	wire source_2_rst;
	wire [1 : 0]source_2_out1_data;
	wire source_2_out1_ready;
	wire source_2_out1_valid;

	wire source_3_clk;
	wire source_3_rst;
	wire [0 : 0]source_3_out1_data;
	wire source_3_out1_ready;
	wire source_3_out1_valid;

	wire source_4_clk;
	wire source_4_rst;
	wire [3 : 0]source_4_out1_data;
	wire source_4_out1_ready;
	wire source_4_out1_valid;

	wire fork_79_clk;
	wire fork_79_rst;
	wire [0 : 0]fork_79_in1_data;
	wire fork_79_in1_ready;
	wire fork_79_in1_valid;
	wire [0 : 0]fork_79_out1_data;
	wire fork_79_out1_ready;
	wire fork_79_out1_valid;
	wire [0 : 0]fork_79_out2_data;
	wire fork_79_out2_ready;
	wire fork_79_out2_valid;

	wire phi_84_clk;
	wire phi_84_rst;
	wire [0 : 0]phi_84_in1_data;
	wire phi_84_in1_ready;
	wire phi_84_in1_valid;
	wire [31 : 0]phi_84_in2_data;
	wire phi_84_in2_ready;
	wire phi_84_in2_valid;
	wire [31 : 0]phi_84_in3_data;
	wire phi_84_in3_ready;
	wire phi_84_in3_valid;
	wire [31 : 0]phi_84_out1_data;
	wire phi_84_out1_ready;
	wire phi_84_out1_valid;

	wire phi_85_clk;
	wire phi_85_rst;
	wire [0 : 0]phi_85_in1_data;
	wire phi_85_in1_ready;
	wire phi_85_in1_valid;
	wire [3 : 0]phi_85_in2_data;
	wire phi_85_in2_ready;
	wire phi_85_in2_valid;
	wire [3 : 0]phi_85_in3_data;
	wire phi_85_in3_ready;
	wire phi_85_in3_valid;
	wire [3 : 0]phi_85_out1_data;
	wire phi_85_out1_ready;
	wire phi_85_out1_valid;

	wire cst_30_clk;
	wire cst_30_rst;
	wire [1 : 0]cst_30_in1_data;
	wire cst_30_in1_ready;
	wire cst_30_in1_valid;
	wire [1 : 0]cst_30_out1_data;
	wire cst_30_out1_ready;
	wire cst_30_out1_valid;

	wire shl_86_clk;
	wire shl_86_rst;
	wire [6 : 0]shl_86_in1_data;
	wire shl_86_in1_ready;
	wire shl_86_in1_valid;
	wire [6 : 0]shl_86_in2_data;
	wire shl_86_in2_ready;
	wire shl_86_in2_valid;
	wire [6 : 0]shl_86_out1_data;
	wire shl_86_out1_ready;
	wire shl_86_out1_valid;

	wire add_87_clk;
	wire add_87_rst;
	wire [7 : 0]add_87_in1_data;
	wire add_87_in1_ready;
	wire add_87_in1_valid;
	wire [7 : 0]add_87_in2_data;
	wire add_87_in2_ready;
	wire add_87_in2_valid;
	wire [7 : 0]add_87_out1_data;
	wire add_87_out1_ready;
	wire add_87_out1_valid;

	wire load_90_clk;
	wire load_90_rst;
	wire [31 : 0]load_90_in1_data;
	wire load_90_in1_ready;
	wire load_90_in1_valid;
	wire [7 : 0]load_90_in2_data;
	wire load_90_in2_ready;
	wire load_90_in2_valid;
	wire [31 : 0]load_90_out1_data;
	wire load_90_out1_ready;
	wire load_90_out1_valid;
	wire [7 : 0]load_90_out2_data;
	wire load_90_out2_ready;
	wire load_90_out2_valid;

	wire cst_31_clk;
	wire cst_31_rst;
	wire [1 : 0]cst_31_in1_data;
	wire cst_31_in1_ready;
	wire cst_31_in1_valid;
	wire [1 : 0]cst_31_out1_data;
	wire cst_31_out1_ready;
	wire cst_31_out1_valid;

	wire shl_91_clk;
	wire shl_91_rst;
	wire [6 : 0]shl_91_in1_data;
	wire shl_91_in1_ready;
	wire shl_91_in1_valid;
	wire [6 : 0]shl_91_in2_data;
	wire shl_91_in2_ready;
	wire shl_91_in2_valid;
	wire [6 : 0]shl_91_out1_data;
	wire shl_91_out1_ready;
	wire shl_91_out1_valid;

	wire add_92_clk;
	wire add_92_rst;
	wire [7 : 0]add_92_in1_data;
	wire add_92_in1_ready;
	wire add_92_in1_valid;
	wire [7 : 0]add_92_in2_data;
	wire add_92_in2_ready;
	wire add_92_in2_valid;
	wire [7 : 0]add_92_out1_data;
	wire add_92_out1_ready;
	wire add_92_out1_valid;

	wire load_95_clk;
	wire load_95_rst;
	wire [31 : 0]load_95_in1_data;
	wire load_95_in1_ready;
	wire load_95_in1_valid;
	wire [7 : 0]load_95_in2_data;
	wire load_95_in2_ready;
	wire load_95_in2_valid;
	wire [31 : 0]load_95_out1_data;
	wire load_95_out1_ready;
	wire load_95_out1_valid;
	wire [7 : 0]load_95_out2_data;
	wire load_95_out2_ready;
	wire load_95_out2_valid;

	wire cst_32_clk;
	wire cst_32_rst;
	wire [0 : 0]cst_32_in1_data;
	wire cst_32_in1_ready;
	wire cst_32_in1_valid;
	wire [0 : 0]cst_32_out1_data;
	wire cst_32_out1_ready;
	wire cst_32_out1_valid;

	wire add_98_clk;
	wire add_98_rst;
	wire [3 : 0]add_98_in1_data;
	wire add_98_in1_ready;
	wire add_98_in1_valid;
	wire [3 : 0]add_98_in2_data;
	wire add_98_in2_ready;
	wire add_98_in2_valid;
	wire [3 : 0]add_98_out1_data;
	wire add_98_out1_ready;
	wire add_98_out1_valid;

	wire cst_33_clk;
	wire cst_33_rst;
	wire [3 : 0]cst_33_in1_data;
	wire cst_33_in1_ready;
	wire cst_33_in1_valid;
	wire [3 : 0]cst_33_out1_data;
	wire cst_33_out1_ready;
	wire cst_33_out1_valid;

	wire icmp_99_clk;
	wire icmp_99_rst;
	wire [3 : 0]icmp_99_in1_data;
	wire icmp_99_in1_ready;
	wire icmp_99_in1_valid;
	wire [3 : 0]icmp_99_in2_data;
	wire icmp_99_in2_ready;
	wire icmp_99_in2_valid;
	wire [0 : 0]icmp_99_out1_data;
	wire icmp_99_out1_ready;
	wire icmp_99_out1_valid;

	wire phi_n19_clk;
	wire phi_n19_rst;
	wire [3 : 0]phi_n19_in1_data;
	wire phi_n19_in1_ready;
	wire phi_n19_in1_valid;
	wire [3 : 0]phi_n19_in2_data;
	wire phi_n19_in2_ready;
	wire phi_n19_in2_valid;
	wire [3 : 0]phi_n19_out1_data;
	wire phi_n19_out1_ready;
	wire phi_n19_out1_valid;

	wire phi_n20_clk;
	wire phi_n20_rst;
	wire [3 : 0]phi_n20_in1_data;
	wire phi_n20_in1_ready;
	wire phi_n20_in1_valid;
	wire [3 : 0]phi_n20_in2_data;
	wire phi_n20_in2_ready;
	wire phi_n20_in2_valid;
	wire [3 : 0]phi_n20_out1_data;
	wire phi_n20_out1_ready;
	wire phi_n20_out1_valid;

	wire fork_13_clk;
	wire fork_13_rst;
	wire [3 : 0]fork_13_in1_data;
	wire fork_13_in1_ready;
	wire fork_13_in1_valid;
	wire [3 : 0]fork_13_out1_data;
	wire fork_13_out1_ready;
	wire fork_13_out1_valid;
	wire [3 : 0]fork_13_out2_data;
	wire fork_13_out2_ready;
	wire fork_13_out2_valid;
	wire [3 : 0]fork_13_out3_data;
	wire fork_13_out3_ready;
	wire fork_13_out3_valid;

	wire fork_15_clk;
	wire fork_15_rst;
	wire [3 : 0]fork_15_in1_data;
	wire fork_15_in1_ready;
	wire fork_15_in1_valid;
	wire [3 : 0]fork_15_out1_data;
	wire fork_15_out1_ready;
	wire fork_15_out1_valid;
	wire [3 : 0]fork_15_out2_data;
	wire fork_15_out2_ready;
	wire fork_15_out2_valid;

	wire fork_31_clk;
	wire fork_31_rst;
	wire [3 : 0]fork_31_in1_data;
	wire fork_31_in1_ready;
	wire fork_31_in1_valid;
	wire [3 : 0]fork_31_out1_data;
	wire fork_31_out1_ready;
	wire fork_31_out1_valid;
	wire [3 : 0]fork_31_out2_data;
	wire fork_31_out2_ready;
	wire fork_31_out2_valid;

	wire fork_32_clk;
	wire fork_32_rst;
	wire [3 : 0]fork_32_in1_data;
	wire fork_32_in1_ready;
	wire fork_32_in1_valid;
	wire [3 : 0]fork_32_out1_data;
	wire fork_32_out1_ready;
	wire fork_32_out1_valid;
	wire [3 : 0]fork_32_out2_data;
	wire fork_32_out2_ready;
	wire fork_32_out2_valid;

	wire branch_35_clk;
	wire branch_35_rst;
	wire [31 : 0]branch_35_in1_data;
	wire branch_35_in1_ready;
	wire branch_35_in1_valid;
	wire [0 : 0]branch_35_in2_data;
	wire branch_35_in2_ready;
	wire branch_35_in2_valid;
	wire [31 : 0]branch_35_out1_data;
	wire branch_35_out1_ready;
	wire branch_35_out1_valid;
	wire [31 : 0]branch_35_out2_data;
	wire branch_35_out2_ready;
	wire branch_35_out2_valid;

	wire branch_36_clk;
	wire branch_36_rst;
	wire [3 : 0]branch_36_in1_data;
	wire branch_36_in1_ready;
	wire branch_36_in1_valid;
	wire [0 : 0]branch_36_in2_data;
	wire branch_36_in2_ready;
	wire branch_36_in2_valid;
	wire [3 : 0]branch_36_out1_data;
	wire branch_36_out1_ready;
	wire branch_36_out1_valid;
	wire [3 : 0]branch_36_out2_data;
	wire branch_36_out2_ready;
	wire branch_36_out2_valid;

	wire branch_37_clk;
	wire branch_37_rst;
	wire [3 : 0]branch_37_in1_data;
	wire branch_37_in1_ready;
	wire branch_37_in1_valid;
	wire [0 : 0]branch_37_in2_data;
	wire branch_37_in2_ready;
	wire branch_37_in2_valid;
	wire [3 : 0]branch_37_out1_data;
	wire branch_37_out1_ready;
	wire branch_37_out1_valid;
	wire [3 : 0]branch_37_out2_data;
	wire branch_37_out2_ready;
	wire branch_37_out2_valid;

	wire branch_38_clk;
	wire branch_38_rst;
	wire [3 : 0]branch_38_in1_data;
	wire branch_38_in1_ready;
	wire branch_38_in1_valid;
	wire [0 : 0]branch_38_in2_data;
	wire branch_38_in2_ready;
	wire branch_38_in2_valid;
	wire [3 : 0]branch_38_out1_data;
	wire branch_38_out1_ready;
	wire branch_38_out1_valid;
	wire [3 : 0]branch_38_out2_data;
	wire branch_38_out2_ready;
	wire branch_38_out2_valid;

	wire fork_48_clk;
	wire fork_48_rst;
	wire [0 : 0]fork_48_in1_data;
	wire fork_48_in1_ready;
	wire fork_48_in1_valid;
	wire [0 : 0]fork_48_out1_data;
	wire fork_48_out1_ready;
	wire fork_48_out1_valid;
	wire [0 : 0]fork_48_out2_data;
	wire fork_48_out2_ready;
	wire fork_48_out2_valid;
	wire [0 : 0]fork_48_out3_data;
	wire fork_48_out3_ready;
	wire fork_48_out3_valid;
	wire [0 : 0]fork_48_out4_data;
	wire fork_48_out4_ready;
	wire fork_48_out4_valid;
	wire [0 : 0]fork_48_out5_data;
	wire fork_48_out5_ready;
	wire fork_48_out5_valid;

	wire phiC_35_clk;
	wire phiC_35_rst;
	wire [0 : 0]phiC_35_in1_data;
	wire phiC_35_in1_ready;
	wire phiC_35_in1_valid;
	wire [0 : 0]phiC_35_in2_data;
	wire phiC_35_in2_ready;
	wire phiC_35_in2_valid;
	wire [0 : 0]phiC_35_out1_data;
	wire phiC_35_out1_ready;
	wire phiC_35_out1_valid;
	wire [0 : 0]phiC_35_out2_data;
	wire phiC_35_out2_ready;
	wire phiC_35_out2_valid;

	wire branchC_57_clk;
	wire branchC_57_rst;
	wire [0 : 0]branchC_57_in1_data;
	wire branchC_57_in1_ready;
	wire branchC_57_in1_valid;
	wire [0 : 0]branchC_57_in2_data;
	wire branchC_57_in2_ready;
	wire branchC_57_in2_valid;
	wire [0 : 0]branchC_57_out1_data;
	wire branchC_57_out1_ready;
	wire branchC_57_out1_valid;
	wire [0 : 0]branchC_57_out2_data;
	wire branchC_57_out2_ready;
	wire branchC_57_out2_valid;

	wire source_21_clk;
	wire source_21_rst;
	wire [1 : 0]source_21_out1_data;
	wire source_21_out1_ready;
	wire source_21_out1_valid;

	wire source_22_clk;
	wire source_22_rst;
	wire [1 : 0]source_22_out1_data;
	wire source_22_out1_ready;
	wire source_22_out1_valid;

	wire source_23_clk;
	wire source_23_rst;
	wire [0 : 0]source_23_out1_data;
	wire source_23_out1_ready;
	wire source_23_out1_valid;

	wire source_24_clk;
	wire source_24_rst;
	wire [3 : 0]source_24_out1_data;
	wire source_24_out1_ready;
	wire source_24_out1_valid;

	wire fork_85_clk;
	wire fork_85_rst;
	wire [0 : 0]fork_85_in1_data;
	wire fork_85_in1_ready;
	wire fork_85_in1_valid;
	wire [0 : 0]fork_85_out1_data;
	wire fork_85_out1_ready;
	wire fork_85_out1_valid;
	wire [0 : 0]fork_85_out2_data;
	wire fork_85_out2_ready;
	wire fork_85_out2_valid;

	wire phi_1_clk;
	wire phi_1_rst;
	wire [0 : 0]phi_1_in1_data;
	wire phi_1_in1_ready;
	wire phi_1_in1_valid;
	wire [3 : 0]phi_1_in2_data;
	wire phi_1_in2_ready;
	wire phi_1_in2_valid;
	wire [3 : 0]phi_1_in3_data;
	wire phi_1_in3_ready;
	wire phi_1_in3_valid;
	wire [3 : 0]phi_1_out1_data;
	wire phi_1_out1_ready;
	wire phi_1_out1_valid;

	wire brCst_block2_clk;
	wire brCst_block2_rst;
	wire [0 : 0]brCst_block2_in1_data;
	wire brCst_block2_in1_ready;
	wire brCst_block2_in1_valid;
	wire [0 : 0]brCst_block2_out1_data;
	wire brCst_block2_out1_ready;
	wire brCst_block2_out1_valid;

	wire cst_1_clk;
	wire cst_1_rst;
	wire [0 : 0]cst_1_in1_data;
	wire cst_1_in1_ready;
	wire cst_1_in1_valid;
	wire [0 : 0]cst_1_out1_data;
	wire cst_1_out1_ready;
	wire cst_1_out1_valid;

	wire branch_1_clk;
	wire branch_1_rst;
	wire [0 : 0]branch_1_in1_data;
	wire branch_1_in1_ready;
	wire branch_1_in1_valid;
	wire [0 : 0]branch_1_in2_data;
	wire branch_1_in2_ready;
	wire branch_1_in2_valid;
	wire [0 : 0]branch_1_out1_data;
	wire branch_1_out1_ready;
	wire branch_1_out1_valid;
	wire [0 : 0]branch_1_out2_data;
	wire branch_1_out2_ready;
	wire branch_1_out2_valid;

	wire branch_2_clk;
	wire branch_2_rst;
	wire [3 : 0]branch_2_in1_data;
	wire branch_2_in1_ready;
	wire branch_2_in1_valid;
	wire [0 : 0]branch_2_in2_data;
	wire branch_2_in2_ready;
	wire branch_2_in2_valid;
	wire [3 : 0]branch_2_out1_data;
	wire branch_2_out1_ready;
	wire branch_2_out1_valid;
	wire [3 : 0]branch_2_out2_data;
	wire branch_2_out2_ready;
	wire branch_2_out2_valid;

	wire fork_34_clk;
	wire fork_34_rst;
	wire [0 : 0]fork_34_in1_data;
	wire fork_34_in1_ready;
	wire fork_34_in1_valid;
	wire [0 : 0]fork_34_out1_data;
	wire fork_34_out1_ready;
	wire fork_34_out1_valid;
	wire [0 : 0]fork_34_out2_data;
	wire fork_34_out2_ready;
	wire fork_34_out2_valid;
	wire [0 : 0]fork_34_out3_data;
	wire fork_34_out3_ready;
	wire fork_34_out3_valid;

	wire phiC_21_clk;
	wire phiC_21_rst;
	wire [0 : 0]phiC_21_in1_data;
	wire phiC_21_in1_ready;
	wire phiC_21_in1_valid;
	wire [0 : 0]phiC_21_in2_data;
	wire phiC_21_in2_ready;
	wire phiC_21_in2_valid;
	wire [0 : 0]phiC_21_out1_data;
	wire phiC_21_out1_ready;
	wire phiC_21_out1_valid;
	wire [0 : 0]phiC_21_out2_data;
	wire phiC_21_out2_ready;
	wire phiC_21_out2_valid;

	wire forkC_54_clk;
	wire forkC_54_rst;
	wire [0 : 0]forkC_54_in1_data;
	wire forkC_54_in1_ready;
	wire forkC_54_in1_valid;
	wire [0 : 0]forkC_54_out1_data;
	wire forkC_54_out1_ready;
	wire forkC_54_out1_valid;
	wire [0 : 0]forkC_54_out2_data;
	wire forkC_54_out2_ready;
	wire forkC_54_out2_valid;
	wire [0 : 0]forkC_54_out3_data;
	wire forkC_54_out3_ready;
	wire forkC_54_out3_valid;

	wire branchC_43_clk;
	wire branchC_43_rst;
	wire [0 : 0]branchC_43_in1_data;
	wire branchC_43_in1_ready;
	wire branchC_43_in1_valid;
	wire [0 : 0]branchC_43_in2_data;
	wire branchC_43_in2_ready;
	wire branchC_43_in2_valid;
	wire [0 : 0]branchC_43_out1_data;
	wire branchC_43_out1_ready;
	wire branchC_43_out1_valid;
	wire [0 : 0]branchC_43_out2_data;
	wire branchC_43_out2_ready;
	wire branchC_43_out2_valid;

	wire MC_E_clk;
	wire MC_E_rst;
	wire [31 : 0]MC_E_in1_data;
	wire MC_E_in1_ready;
	wire MC_E_in1_valid;
	wire [7 : 0]MC_E_in2_data;
	wire MC_E_in2_ready;
	wire MC_E_in2_valid;
	wire [7 : 0]MC_E_in3_data;
	wire MC_E_in3_ready;
	wire MC_E_in3_valid;
	wire [31 : 0]MC_E_in4_data;
	wire MC_E_in4_ready;
	wire MC_E_in4_valid;
	wire [7 : 0]MC_E_in5_data;
	wire MC_E_in5_ready;
	wire MC_E_in5_valid;
	wire [31 : 0]MC_E_out1_data;
	wire MC_E_out1_ready;
	wire MC_E_out1_valid;
	wire [31 : 0]MC_E_out2_data;
	wire MC_E_out2_ready;
	wire MC_E_out2_valid;
	wire [0 : 0]MC_E_out3_data;
	wire MC_E_out3_ready;
	wire MC_E_out3_valid;

	wire MC_A_clk;
	wire MC_A_rst;
	wire [7 : 0]MC_A_in1_data;
	wire MC_A_in1_ready;
	wire MC_A_in1_valid;
	wire [31 : 0]MC_A_in2_data;
	wire MC_A_in2_ready;
	wire MC_A_in2_valid;
	wire [7 : 0]MC_A_in3_data;
	wire MC_A_in3_ready;
	wire MC_A_in3_valid;
	wire [31 : 0]MC_A_in4_data;
	wire MC_A_in4_ready;
	wire MC_A_in4_valid;
	wire [31 : 0]MC_A_out1_data;
	wire MC_A_out1_ready;
	wire MC_A_out1_valid;
	wire [0 : 0]MC_A_out2_data;
	wire MC_A_out2_ready;
	wire MC_A_out2_valid;

	wire MC_B_clk;
	wire MC_B_rst;
	wire [7 : 0]MC_B_in1_data;
	wire MC_B_in1_ready;
	wire MC_B_in1_valid;
	wire [31 : 0]MC_B_in2_data;
	wire MC_B_in2_ready;
	wire MC_B_in2_valid;
	wire [7 : 0]MC_B_in3_data;
	wire MC_B_in3_ready;
	wire MC_B_in3_valid;
	wire [31 : 0]MC_B_in4_data;
	wire MC_B_in4_ready;
	wire MC_B_in4_valid;
	wire [31 : 0]MC_B_out1_data;
	wire MC_B_out1_ready;
	wire MC_B_out1_valid;
	wire [0 : 0]MC_B_out2_data;
	wire MC_B_out2_ready;
	wire MC_B_out2_valid;

	wire MC_F_clk;
	wire MC_F_rst;
	wire [31 : 0]MC_F_in1_data;
	wire MC_F_in1_ready;
	wire MC_F_in1_valid;
	wire [7 : 0]MC_F_in2_data;
	wire MC_F_in2_ready;
	wire MC_F_in2_valid;
	wire [7 : 0]MC_F_in3_data;
	wire MC_F_in3_ready;
	wire MC_F_in3_valid;
	wire [31 : 0]MC_F_in4_data;
	wire MC_F_in4_ready;
	wire MC_F_in4_valid;
	wire [7 : 0]MC_F_in5_data;
	wire MC_F_in5_ready;
	wire MC_F_in5_valid;
	wire [31 : 0]MC_F_out1_data;
	wire MC_F_out1_ready;
	wire MC_F_out1_valid;
	wire [31 : 0]MC_F_out2_data;
	wire MC_F_out2_ready;
	wire MC_F_out2_valid;
	wire [0 : 0]MC_F_out3_data;
	wire MC_F_out3_ready;
	wire MC_F_out3_valid;

	wire MC_C_clk;
	wire MC_C_rst;
	wire [7 : 0]MC_C_in1_data;
	wire MC_C_in1_ready;
	wire MC_C_in1_valid;
	wire [31 : 0]MC_C_in2_data;
	wire MC_C_in2_ready;
	wire MC_C_in2_valid;
	wire [7 : 0]MC_C_in3_data;
	wire MC_C_in3_ready;
	wire MC_C_in3_valid;
	wire [31 : 0]MC_C_in4_data;
	wire MC_C_in4_ready;
	wire MC_C_in4_valid;
	wire [31 : 0]MC_C_out1_data;
	wire MC_C_out1_ready;
	wire MC_C_out1_valid;
	wire [0 : 0]MC_C_out2_data;
	wire MC_C_out2_ready;
	wire MC_C_out2_valid;

	wire MC_D_clk;
	wire MC_D_rst;
	wire [7 : 0]MC_D_in1_data;
	wire MC_D_in1_ready;
	wire MC_D_in1_valid;
	wire [31 : 0]MC_D_in2_data;
	wire MC_D_in2_ready;
	wire MC_D_in2_valid;
	wire [7 : 0]MC_D_in3_data;
	wire MC_D_in3_ready;
	wire MC_D_in3_valid;
	wire [31 : 0]MC_D_in4_data;
	wire MC_D_in4_ready;
	wire MC_D_in4_valid;
	wire [31 : 0]MC_D_out1_data;
	wire MC_D_out1_ready;
	wire MC_D_out1_valid;
	wire [0 : 0]MC_D_out2_data;
	wire MC_D_out2_ready;
	wire MC_D_out2_valid;

	wire MC_G_clk;
	wire MC_G_rst;
	wire [31 : 0]MC_G_in1_data;
	wire MC_G_in1_ready;
	wire MC_G_in1_valid;
	wire [7 : 0]MC_G_in2_data;
	wire MC_G_in2_ready;
	wire MC_G_in2_valid;
	wire [7 : 0]MC_G_in3_data;
	wire MC_G_in3_ready;
	wire MC_G_in3_valid;
	wire [31 : 0]MC_G_in4_data;
	wire MC_G_in4_ready;
	wire MC_G_in4_valid;
	wire [31 : 0]MC_G_out1_data;
	wire MC_G_out1_ready;
	wire MC_G_out1_valid;
	wire [0 : 0]MC_G_out2_data;
	wire MC_G_out2_ready;
	wire MC_G_out2_valid;

	wire sink_0_clk;
	wire sink_0_rst;
	wire [0 : 0]sink_0_in1_data;
	wire sink_0_in1_ready;
	wire sink_0_in1_valid;

	wire sink_1_clk;
	wire sink_1_rst;
	wire [0 : 0]sink_1_in1_data;
	wire sink_1_in1_ready;
	wire sink_1_in1_valid;

	wire sink_2_clk;
	wire sink_2_rst;
	wire [3 : 0]sink_2_in1_data;
	wire sink_2_in1_ready;
	wire sink_2_in1_valid;

	wire sink_3_clk;
	wire sink_3_rst;
	wire [31 : 0]sink_3_in1_data;
	wire sink_3_in1_ready;
	wire sink_3_in1_valid;

	wire sink_4_clk;
	wire sink_4_rst;
	wire [0 : 0]sink_4_in1_data;
	wire sink_4_in1_ready;
	wire sink_4_in1_valid;

	wire sink_5_clk;
	wire sink_5_rst;
	wire [3 : 0]sink_5_in1_data;
	wire sink_5_in1_ready;
	wire sink_5_in1_valid;

	wire sink_6_clk;
	wire sink_6_rst;
	wire [3 : 0]sink_6_in1_data;
	wire sink_6_in1_ready;
	wire sink_6_in1_valid;

	wire sink_7_clk;
	wire sink_7_rst;
	wire [3 : 0]sink_7_in1_data;
	wire sink_7_in1_ready;
	wire sink_7_in1_valid;

	wire sink_8_clk;
	wire sink_8_rst;
	wire [3 : 0]sink_8_in1_data;
	wire sink_8_in1_ready;
	wire sink_8_in1_valid;

	wire sink_9_clk;
	wire sink_9_rst;
	wire [3 : 0]sink_9_in1_data;
	wire sink_9_in1_ready;
	wire sink_9_in1_valid;

	wire sink_10_clk;
	wire sink_10_rst;
	wire [0 : 0]sink_10_in1_data;
	wire sink_10_in1_ready;
	wire sink_10_in1_valid;

	wire sink_11_clk;
	wire sink_11_rst;
	wire [0 : 0]sink_11_in1_data;
	wire sink_11_in1_ready;
	wire sink_11_in1_valid;

	wire sink_12_clk;
	wire sink_12_rst;
	wire [3 : 0]sink_12_in1_data;
	wire sink_12_in1_ready;
	wire sink_12_in1_valid;

	wire sink_13_clk;
	wire sink_13_rst;
	wire [31 : 0]sink_13_in1_data;
	wire sink_13_in1_ready;
	wire sink_13_in1_valid;

	wire sink_14_clk;
	wire sink_14_rst;
	wire [0 : 0]sink_14_in1_data;
	wire sink_14_in1_ready;
	wire sink_14_in1_valid;

	wire sink_15_clk;
	wire sink_15_rst;
	wire [3 : 0]sink_15_in1_data;
	wire sink_15_in1_ready;
	wire sink_15_in1_valid;

	wire sink_16_clk;
	wire sink_16_rst;
	wire [3 : 0]sink_16_in1_data;
	wire sink_16_in1_ready;
	wire sink_16_in1_valid;

	wire sink_17_clk;
	wire sink_17_rst;
	wire [3 : 0]sink_17_in1_data;
	wire sink_17_in1_ready;
	wire sink_17_in1_valid;

	wire sink_18_clk;
	wire sink_18_rst;
	wire [3 : 0]sink_18_in1_data;
	wire sink_18_in1_ready;
	wire sink_18_in1_valid;

	wire sink_19_clk;
	wire sink_19_rst;
	wire [3 : 0]sink_19_in1_data;
	wire sink_19_in1_ready;
	wire sink_19_in1_valid;

	wire sink_20_clk;
	wire sink_20_rst;
	wire [0 : 0]sink_20_in1_data;
	wire sink_20_in1_ready;
	wire sink_20_in1_valid;

	wire sink_21_clk;
	wire sink_21_rst;
	wire [0 : 0]sink_21_in1_data;
	wire sink_21_in1_ready;
	wire sink_21_in1_valid;

	wire sink_22_clk;
	wire sink_22_rst;
	wire [3 : 0]sink_22_in1_data;
	wire sink_22_in1_ready;
	wire sink_22_in1_valid;

	wire sink_23_clk;
	wire sink_23_rst;
	wire [31 : 0]sink_23_in1_data;
	wire sink_23_in1_ready;
	wire sink_23_in1_valid;

	wire sink_24_clk;
	wire sink_24_rst;
	wire [0 : 0]sink_24_in1_data;
	wire sink_24_in1_ready;
	wire sink_24_in1_valid;

	wire sink_25_clk;
	wire sink_25_rst;
	wire [3 : 0]sink_25_in1_data;
	wire sink_25_in1_ready;
	wire sink_25_in1_valid;

	wire sink_26_clk;
	wire sink_26_rst;
	wire [3 : 0]sink_26_in1_data;
	wire sink_26_in1_ready;
	wire sink_26_in1_valid;

	wire sink_27_clk;
	wire sink_27_rst;
	wire [3 : 0]sink_27_in1_data;
	wire sink_27_in1_ready;
	wire sink_27_in1_valid;

	wire sink_28_clk;
	wire sink_28_rst;
	wire [3 : 0]sink_28_in1_data;
	wire sink_28_in1_ready;
	wire sink_28_in1_valid;

	wire sink_29_clk;
	wire sink_29_rst;
	wire [3 : 0]sink_29_in1_data;
	wire sink_29_in1_ready;
	wire sink_29_in1_valid;

	wire sink_30_clk;
	wire sink_30_rst;
	wire [0 : 0]sink_30_in1_data;
	wire sink_30_in1_ready;
	wire sink_30_in1_valid;

	wire sink_31_clk;
	wire sink_31_rst;
	wire [0 : 0]sink_31_in1_data;
	wire sink_31_in1_ready;
	wire sink_31_in1_valid;

	wire sink_32_clk;
	wire sink_32_rst;
	wire [0 : 0]sink_32_in1_data;
	wire sink_32_in1_ready;
	wire sink_32_in1_valid;

	wire sink_33_clk;
	wire sink_33_rst;
	wire [0 : 0]sink_33_in1_data;
	wire sink_33_in1_ready;
	wire sink_33_in1_valid;

	wire sink_34_clk;
	wire sink_34_rst;
	wire [0 : 0]sink_34_in1_data;
	wire sink_34_in1_ready;
	wire sink_34_in1_valid;

	wire sink_35_clk;
	wire sink_35_rst;
	wire [0 : 0]sink_35_in1_data;
	wire sink_35_in1_ready;
	wire sink_35_in1_valid;

	wire sink_36_clk;
	wire sink_36_rst;
	wire [0 : 0]sink_36_in1_data;
	wire sink_36_in1_ready;
	wire sink_36_in1_valid;

	wire sink_37_clk;
	wire sink_37_rst;
	wire [0 : 0]sink_37_in1_data;
	wire sink_37_in1_ready;
	wire sink_37_in1_valid;

	wire sink_38_clk;
	wire sink_38_rst;
	wire [0 : 0]sink_38_in1_data;
	wire sink_38_in1_ready;
	wire sink_38_in1_valid;

	wire Buffer_100_clk;
	wire Buffer_100_rst;
	wire [31 : 0]Buffer_100_in1_data;
	wire Buffer_100_in1_ready;
	wire Buffer_100_in1_valid;
	wire [31 : 0]Buffer_100_out1_data;
	wire Buffer_100_out1_ready;
	wire Buffer_100_out1_valid;

	wire Buffer_101_clk;
	wire Buffer_101_rst;
	wire [31 : 0]Buffer_101_in1_data;
	wire Buffer_101_in1_ready;
	wire Buffer_101_in1_valid;
	wire [31 : 0]Buffer_101_out1_data;
	wire Buffer_101_out1_ready;
	wire Buffer_101_out1_valid;

	wire Buffer_102_clk;
	wire Buffer_102_rst;
	wire [31 : 0]Buffer_102_in1_data;
	wire Buffer_102_in1_ready;
	wire Buffer_102_in1_valid;
	wire [31 : 0]Buffer_102_out1_data;
	wire Buffer_102_out1_ready;
	wire Buffer_102_out1_valid;

	wire Buffer_103_clk;
	wire Buffer_103_rst;
	wire [31 : 0]Buffer_103_in1_data;
	wire Buffer_103_in1_ready;
	wire Buffer_103_in1_valid;
	wire [31 : 0]Buffer_103_out1_data;
	wire Buffer_103_out1_ready;
	wire Buffer_103_out1_valid;

	wire Buffer_104_clk;
	wire Buffer_104_rst;
	wire [31 : 0]Buffer_104_in1_data;
	wire Buffer_104_in1_ready;
	wire Buffer_104_in1_valid;
	wire [31 : 0]Buffer_104_out1_data;
	wire Buffer_104_out1_ready;
	wire Buffer_104_out1_valid;

	wire Buffer_105_clk;
	wire Buffer_105_rst;
	wire [31 : 0]Buffer_105_in1_data;
	wire Buffer_105_in1_ready;
	wire Buffer_105_in1_valid;
	wire [31 : 0]Buffer_105_out1_data;
	wire Buffer_105_out1_ready;
	wire Buffer_105_out1_valid;

	wire Buffer_106_clk;
	wire Buffer_106_rst;
	wire [31 : 0]Buffer_106_in1_data;
	wire Buffer_106_in1_ready;
	wire Buffer_106_in1_valid;
	wire [31 : 0]Buffer_106_out1_data;
	wire Buffer_106_out1_ready;
	wire Buffer_106_out1_valid;

	wire Buffer_107_clk;
	wire Buffer_107_rst;
	wire [31 : 0]Buffer_107_in1_data;
	wire Buffer_107_in1_ready;
	wire Buffer_107_in1_valid;
	wire [31 : 0]Buffer_107_out1_data;
	wire Buffer_107_out1_ready;
	wire Buffer_107_out1_valid;

	wire Buffer_108_clk;
	wire Buffer_108_rst;
	wire [31 : 0]Buffer_108_in1_data;
	wire Buffer_108_in1_ready;
	wire Buffer_108_in1_valid;
	wire [31 : 0]Buffer_108_out1_data;
	wire Buffer_108_out1_ready;
	wire Buffer_108_out1_valid;

	wire Buffer_109_clk;
	wire Buffer_109_rst;
	wire [31 : 0]Buffer_109_in1_data;
	wire Buffer_109_in1_ready;
	wire Buffer_109_in1_valid;
	wire [31 : 0]Buffer_109_out1_data;
	wire Buffer_109_out1_ready;
	wire Buffer_109_out1_valid;

	wire Buffer_110_clk;
	wire Buffer_110_rst;
	wire [31 : 0]Buffer_110_in1_data;
	wire Buffer_110_in1_ready;
	wire Buffer_110_in1_valid;
	wire [31 : 0]Buffer_110_out1_data;
	wire Buffer_110_out1_ready;
	wire Buffer_110_out1_valid;

	wire Buffer_111_clk;
	wire Buffer_111_rst;
	wire [31 : 0]Buffer_111_in1_data;
	wire Buffer_111_in1_ready;
	wire Buffer_111_in1_valid;
	wire [31 : 0]Buffer_111_out1_data;
	wire Buffer_111_out1_ready;
	wire Buffer_111_out1_valid;

	wire Buffer_112_clk;
	wire Buffer_112_rst;
	wire [31 : 0]Buffer_112_in1_data;
	wire Buffer_112_in1_ready;
	wire Buffer_112_in1_valid;
	wire [31 : 0]Buffer_112_out1_data;
	wire Buffer_112_out1_ready;
	wire Buffer_112_out1_valid;

	wire Buffer_113_clk;
	wire Buffer_113_rst;
	wire [31 : 0]Buffer_113_in1_data;
	wire Buffer_113_in1_ready;
	wire Buffer_113_in1_valid;
	wire [31 : 0]Buffer_113_out1_data;
	wire Buffer_113_out1_ready;
	wire Buffer_113_out1_valid;

	wire Buffer_114_clk;
	wire Buffer_114_rst;
	wire [31 : 0]Buffer_114_in1_data;
	wire Buffer_114_in1_ready;
	wire Buffer_114_in1_valid;
	wire [31 : 0]Buffer_114_out1_data;
	wire Buffer_114_out1_ready;
	wire Buffer_114_out1_valid;

	wire Buffer_115_clk;
	wire Buffer_115_rst;
	wire [31 : 0]Buffer_115_in1_data;
	wire Buffer_115_in1_ready;
	wire Buffer_115_in1_valid;
	wire [31 : 0]Buffer_115_out1_data;
	wire Buffer_115_out1_ready;
	wire Buffer_115_out1_valid;

	wire Buffer_116_clk;
	wire Buffer_116_rst;
	wire [31 : 0]Buffer_116_in1_data;
	wire Buffer_116_in1_ready;
	wire Buffer_116_in1_valid;
	wire [31 : 0]Buffer_116_out1_data;
	wire Buffer_116_out1_ready;
	wire Buffer_116_out1_valid;

	wire Buffer_117_clk;
	wire Buffer_117_rst;
	wire [31 : 0]Buffer_117_in1_data;
	wire Buffer_117_in1_ready;
	wire Buffer_117_in1_valid;
	wire [31 : 0]Buffer_117_out1_data;
	wire Buffer_117_out1_ready;
	wire Buffer_117_out1_valid;

	wire Buffer_118_clk;
	wire Buffer_118_rst;
	wire [31 : 0]Buffer_118_in1_data;
	wire Buffer_118_in1_ready;
	wire Buffer_118_in1_valid;
	wire [31 : 0]Buffer_118_out1_data;
	wire Buffer_118_out1_ready;
	wire Buffer_118_out1_valid;

	wire Buffer_119_clk;
	wire Buffer_119_rst;
	wire [31 : 0]Buffer_119_in1_data;
	wire Buffer_119_in1_ready;
	wire Buffer_119_in1_valid;
	wire [31 : 0]Buffer_119_out1_data;
	wire Buffer_119_out1_ready;
	wire Buffer_119_out1_valid;

	wire Buffer_120_clk;
	wire Buffer_120_rst;
	wire [31 : 0]Buffer_120_in1_data;
	wire Buffer_120_in1_ready;
	wire Buffer_120_in1_valid;
	wire [31 : 0]Buffer_120_out1_data;
	wire Buffer_120_out1_ready;
	wire Buffer_120_out1_valid;

	wire Buffer_121_clk;
	wire Buffer_121_rst;
	wire [31 : 0]Buffer_121_in1_data;
	wire Buffer_121_in1_ready;
	wire Buffer_121_in1_valid;
	wire [31 : 0]Buffer_121_out1_data;
	wire Buffer_121_out1_ready;
	wire Buffer_121_out1_valid;

	wire Buffer_122_clk;
	wire Buffer_122_rst;
	wire [31 : 0]Buffer_122_in1_data;
	wire Buffer_122_in1_ready;
	wire Buffer_122_in1_valid;
	wire [31 : 0]Buffer_122_out1_data;
	wire Buffer_122_out1_ready;
	wire Buffer_122_out1_valid;

	wire Buffer_123_clk;
	wire Buffer_123_rst;
	wire [31 : 0]Buffer_123_in1_data;
	wire Buffer_123_in1_ready;
	wire Buffer_123_in1_valid;
	wire [31 : 0]Buffer_123_out1_data;
	wire Buffer_123_out1_ready;
	wire Buffer_123_out1_valid;

	wire Buffer_124_clk;
	wire Buffer_124_rst;
	wire [31 : 0]Buffer_124_in1_data;
	wire Buffer_124_in1_ready;
	wire Buffer_124_in1_valid;
	wire [31 : 0]Buffer_124_out1_data;
	wire Buffer_124_out1_ready;
	wire Buffer_124_out1_valid;

	wire Buffer_125_clk;
	wire Buffer_125_rst;
	wire [31 : 0]Buffer_125_in1_data;
	wire Buffer_125_in1_ready;
	wire Buffer_125_in1_valid;
	wire [31 : 0]Buffer_125_out1_data;
	wire Buffer_125_out1_ready;
	wire Buffer_125_out1_valid;

	wire Buffer_126_clk;
	wire Buffer_126_rst;
	wire [31 : 0]Buffer_126_in1_data;
	wire Buffer_126_in1_ready;
	wire Buffer_126_in1_valid;
	wire [31 : 0]Buffer_126_out1_data;
	wire Buffer_126_out1_ready;
	wire Buffer_126_out1_valid;

	wire Buffer_127_clk;
	wire Buffer_127_rst;
	wire [31 : 0]Buffer_127_in1_data;
	wire Buffer_127_in1_ready;
	wire Buffer_127_in1_valid;
	wire [31 : 0]Buffer_127_out1_data;
	wire Buffer_127_out1_ready;
	wire Buffer_127_out1_valid;

	wire Buffer_128_clk;
	wire Buffer_128_rst;
	wire [31 : 0]Buffer_128_in1_data;
	wire Buffer_128_in1_ready;
	wire Buffer_128_in1_valid;
	wire [31 : 0]Buffer_128_out1_data;
	wire Buffer_128_out1_ready;
	wire Buffer_128_out1_valid;

	wire Buffer_129_clk;
	wire Buffer_129_rst;
	wire [31 : 0]Buffer_129_in1_data;
	wire Buffer_129_in1_ready;
	wire Buffer_129_in1_valid;
	wire [31 : 0]Buffer_129_out1_data;
	wire Buffer_129_out1_ready;
	wire Buffer_129_out1_valid;

	wire and_300_clk;
	wire and_300_rst;
	wire [31 : 0]and_300_in1_data;
	wire and_300_in1_ready;
	wire and_300_in1_valid;
	wire [31 : 0]and_300_in2_data;
	wire and_300_in2_ready;
	wire and_300_in2_valid;
	wire [31 : 0]and_300_out1_data;
	wire and_300_out1_ready;
	wire and_300_out1_valid;

	wire Buffer_300_clk;
	wire Buffer_300_rst;
	wire [31 : 0]Buffer_300_in1_data;
	wire Buffer_300_in1_ready;
	wire Buffer_300_in1_valid;
	wire [31 : 0]Buffer_300_out1_data;
	wire Buffer_300_out1_ready;
	wire Buffer_300_out1_valid;

	wire and_301_clk;
	wire and_301_rst;
	wire [31 : 0]and_301_in1_data;
	wire and_301_in1_ready;
	wire and_301_in1_valid;
	wire [31 : 0]and_301_in2_data;
	wire and_301_in2_ready;
	wire and_301_in2_valid;
	wire [31 : 0]and_301_out1_data;
	wire and_301_out1_ready;
	wire and_301_out1_valid;

	wire Buffer_301_clk;
	wire Buffer_301_rst;
	wire [31 : 0]Buffer_301_in1_data;
	wire Buffer_301_in1_ready;
	wire Buffer_301_in1_valid;
	wire [31 : 0]Buffer_301_out1_data;
	wire Buffer_301_out1_ready;
	wire Buffer_301_out1_valid;

	wire and_302_clk;
	wire and_302_rst;
	wire [31 : 0]and_302_in1_data;
	wire and_302_in1_ready;
	wire and_302_in1_valid;
	wire [31 : 0]and_302_in2_data;
	wire and_302_in2_ready;
	wire and_302_in2_valid;
	wire [31 : 0]and_302_out1_data;
	wire and_302_out1_ready;
	wire and_302_out1_valid;

	wire Buffer_302_clk;
	wire Buffer_302_rst;
	wire [31 : 0]Buffer_302_in1_data;
	wire Buffer_302_in1_ready;
	wire Buffer_302_in1_valid;
	wire [31 : 0]Buffer_302_out1_data;
	wire Buffer_302_out1_ready;
	wire Buffer_302_out1_valid;

	wire and_303_clk;
	wire and_303_rst;
	wire [31 : 0]and_303_in1_data;
	wire and_303_in1_ready;
	wire and_303_in1_valid;
	wire [31 : 0]and_303_in2_data;
	wire and_303_in2_ready;
	wire and_303_in2_valid;
	wire [31 : 0]and_303_out1_data;
	wire and_303_out1_ready;
	wire and_303_out1_valid;

	wire Buffer_303_clk;
	wire Buffer_303_rst;
	wire [31 : 0]Buffer_303_in1_data;
	wire Buffer_303_in1_ready;
	wire Buffer_303_in1_valid;
	wire [31 : 0]Buffer_303_out1_data;
	wire Buffer_303_out1_ready;
	wire Buffer_303_out1_valid;

	wire and_304_clk;
	wire and_304_rst;
	wire [31 : 0]and_304_in1_data;
	wire and_304_in1_ready;
	wire and_304_in1_valid;
	wire [31 : 0]and_304_in2_data;
	wire and_304_in2_ready;
	wire and_304_in2_valid;
	wire [31 : 0]and_304_out1_data;
	wire and_304_out1_ready;
	wire and_304_out1_valid;

	wire Buffer_304_clk;
	wire Buffer_304_rst;
	wire [31 : 0]Buffer_304_in1_data;
	wire Buffer_304_in1_ready;
	wire Buffer_304_in1_valid;
	wire [31 : 0]Buffer_304_out1_data;
	wire Buffer_304_out1_ready;
	wire Buffer_304_out1_valid;

	wire and_305_clk;
	wire and_305_rst;
	wire [31 : 0]and_305_in1_data;
	wire and_305_in1_ready;
	wire and_305_in1_valid;
	wire [31 : 0]and_305_in2_data;
	wire and_305_in2_ready;
	wire and_305_in2_valid;
	wire [31 : 0]and_305_out1_data;
	wire and_305_out1_ready;
	wire and_305_out1_valid;

	wire Buffer_305_clk;
	wire Buffer_305_rst;
	wire [31 : 0]Buffer_305_in1_data;
	wire Buffer_305_in1_ready;
	wire Buffer_305_in1_valid;
	wire [31 : 0]Buffer_305_out1_data;
	wire Buffer_305_out1_ready;
	wire Buffer_305_out1_valid;



	assign phi_3_clk = clk;
	assign phi_3_rst = rst;
	assign fork_0_in1_data = phi_3_out1_data;
	assign fork_0_in1_valid = phi_3_out1_valid;
	assign phi_3_out1_ready = fork_0_in1_ready;

	assign cst_2_clk = clk;
	assign cst_2_rst = rst;
	assign shl_4_in2_data = cst_2_out1_data;
	assign shl_4_in2_valid = cst_2_out1_valid;
	assign cst_2_out1_ready = shl_4_in2_ready;

	assign shl_4_clk = clk;
	assign shl_4_rst = rst;
	assign add_5_in1_data = shl_4_out1_data;
	assign add_5_in1_valid = shl_4_out1_valid;
	assign shl_4_out1_ready = add_5_in1_ready;

	assign add_5_clk = clk;
	assign add_5_rst = rst;
	assign load_8_in2_data = add_5_out1_data;
	assign load_8_in2_valid = add_5_out1_valid;
	assign add_5_out1_ready = load_8_in2_ready;

	assign load_8_clk = clk;
	assign load_8_rst = rst;
	assign branch_3_in1_data = load_8_out1_data;
	assign branch_3_in1_valid = load_8_out1_valid;
	assign load_8_out1_ready = branch_3_in1_ready;
	assign MC_E_in2_data = load_8_out2_data;
	assign MC_E_in2_valid = load_8_out2_valid;
	assign load_8_out2_ready = MC_E_in2_ready;

	assign brCst_block3_clk = clk;
	assign brCst_block3_rst = rst;
	assign fork_35_in1_data = brCst_block3_out1_data;
	assign fork_35_in1_valid = brCst_block3_out1_valid;
	assign brCst_block3_out1_ready = fork_35_in1_ready;

	assign cst_3_clk = clk;
	assign cst_3_rst = rst;
	assign branch_4_in1_data = cst_3_out1_data;
	assign branch_4_in1_valid = cst_3_out1_valid;
	assign cst_3_out1_ready = branch_4_in1_ready;

	assign phi_n4_clk = clk;
	assign phi_n4_rst = rst;
	assign fork_20_in1_data = phi_n4_out1_data;
	assign fork_20_in1_valid = phi_n4_out1_valid;
	assign phi_n4_out1_ready = fork_20_in1_ready;

	assign fork_0_clk = clk;
	assign fork_0_rst = rst;
	assign add_5_in2_data = fork_0_out1_data;
	assign add_5_in2_valid = fork_0_out1_valid;
	assign fork_0_out1_ready = add_5_in2_ready;
	assign branch_5_in1_data = fork_0_out2_data;
	assign branch_5_in1_valid = fork_0_out2_valid;
	assign fork_0_out2_ready = branch_5_in1_ready;

	assign fork_20_clk = clk;
	assign fork_20_rst = rst;
	assign shl_4_in1_data = fork_20_out1_data;
	assign shl_4_in1_valid = fork_20_out1_valid;
	assign fork_20_out1_ready = shl_4_in1_ready;
	assign branch_6_in1_data = fork_20_out2_data;
	assign branch_6_in1_valid = fork_20_out2_valid;
	assign fork_20_out2_ready = branch_6_in1_ready;

	assign branch_3_clk = clk;
	assign branch_3_rst = rst;
	assign phi_10_in2_data = branch_3_out1_data;
	assign phi_10_in2_valid = branch_3_out1_valid;
	assign branch_3_out1_ready = phi_10_in2_ready;
	assign sink_3_in1_data = branch_3_out2_data;
	assign sink_3_in1_valid = branch_3_out2_valid;
	assign branch_3_out2_ready = sink_3_in1_ready;

	assign branch_4_clk = clk;
	assign branch_4_rst = rst;
	assign phi_11_in2_data = branch_4_out1_data;
	assign phi_11_in2_valid = branch_4_out1_valid;
	assign branch_4_out1_ready = phi_11_in2_ready;
	assign sink_4_in1_data = branch_4_out2_data;
	assign sink_4_in1_valid = branch_4_out2_valid;
	assign branch_4_out2_ready = sink_4_in1_ready;

	assign branch_5_clk = clk;
	assign branch_5_rst = rst;
	assign phi_n9_in1_data = branch_5_out1_data;
	assign phi_n9_in1_valid = branch_5_out1_valid;
	assign branch_5_out1_ready = phi_n9_in1_ready;
	assign sink_5_in1_data = branch_5_out2_data;
	assign sink_5_in1_valid = branch_5_out2_valid;
	assign branch_5_out2_ready = sink_5_in1_ready;

	assign branch_6_clk = clk;
	assign branch_6_rst = rst;
	assign phi_n8_in1_data = branch_6_out1_data;
	assign phi_n8_in1_valid = branch_6_out1_valid;
	assign branch_6_out1_ready = phi_n8_in1_ready;
	assign sink_6_in1_data = branch_6_out2_data;
	assign sink_6_in1_valid = branch_6_out2_valid;
	assign branch_6_out2_ready = sink_6_in1_ready;

	assign fork_35_clk = clk;
	assign fork_35_rst = rst;
	assign branch_6_in2_data = fork_35_out1_data;
	assign branch_6_in2_valid = fork_35_out1_valid;
	assign fork_35_out1_ready = branch_6_in2_ready;
	assign branch_5_in2_data = fork_35_out2_data;
	assign branch_5_in2_valid = fork_35_out2_valid;
	assign fork_35_out2_ready = branch_5_in2_ready;
	assign branch_4_in2_data = fork_35_out3_data;
	assign branch_4_in2_valid = fork_35_out3_valid;
	assign fork_35_out3_ready = branch_4_in2_ready;
	assign branch_3_in2_data = fork_35_out4_data;
	assign branch_3_in2_valid = fork_35_out4_valid;
	assign fork_35_out4_ready = branch_3_in2_ready;
	assign branchC_44_in2_data = fork_35_out5_data;
	assign branchC_44_in2_valid = fork_35_out5_valid;
	assign fork_35_out5_ready = branchC_44_in2_ready;

	assign phiC_22_clk = clk;
	assign phiC_22_rst = rst;
	assign forkC_55_in1_data = phiC_22_out1_data;
	assign forkC_55_in1_valid = phiC_22_out1_valid;
	assign phiC_22_out1_ready = forkC_55_in1_ready;
	assign phi_3_in1_data = phiC_22_out2_data;
	assign phi_3_in1_valid = phiC_22_out2_valid;
	assign phiC_22_out2_ready = phi_3_in1_ready;

	assign forkC_55_clk = clk;
	assign forkC_55_rst = rst;
	assign cst_3_in1_data = forkC_55_out1_data;
	assign cst_3_in1_valid = forkC_55_out1_valid;
	assign forkC_55_out1_ready = cst_3_in1_ready;
	assign branchC_44_in1_data = forkC_55_out2_data;
	assign branchC_44_in1_valid = forkC_55_out2_valid;
	assign forkC_55_out2_ready = branchC_44_in1_ready;
	assign brCst_block3_in1_data = forkC_55_out3_data;
	assign brCst_block3_in1_valid = forkC_55_out3_valid;
	assign forkC_55_out3_ready = brCst_block3_in1_ready;

	assign branchC_44_clk = clk;
	assign branchC_44_rst = rst;
	assign phiC_23_in1_data = branchC_44_out1_data;
	assign phiC_23_in1_valid = branchC_44_out1_valid;
	assign branchC_44_out1_ready = phiC_23_in1_ready;
	assign sink_32_in1_data = branchC_44_out2_data;
	assign sink_32_in1_valid = branchC_44_out2_valid;
	assign branchC_44_out2_ready = sink_32_in1_ready;

	assign source_0_clk = clk;
	assign source_0_rst = rst;
	assign cst_2_in1_data = source_0_out1_data;
	assign cst_2_in1_valid = source_0_out1_valid;
	assign source_0_out1_ready = cst_2_in1_ready;

	assign cst_8_clk = clk;
	assign cst_8_rst = rst;
	assign shl_27_in2_data = cst_8_out1_data;
	assign shl_27_in2_valid = cst_8_out1_valid;
	assign cst_8_out1_ready = shl_27_in2_ready;

	assign shl_27_clk = clk;
	assign shl_27_rst = rst;
	assign add_28_in1_data = shl_27_out1_data;
	assign add_28_in1_valid = shl_27_out1_valid;
	assign shl_27_out1_ready = add_28_in1_ready;

	assign add_28_clk = clk;
	assign add_28_rst = rst;
	assign store_0_in2_data = add_28_out1_data;
	assign store_0_in2_valid = add_28_out1_valid;
	assign add_28_out1_ready = store_0_in2_ready;

	assign store_0_clk = clk;
	assign store_0_rst = rst;
	assign MC_E_in4_data = store_0_out1_data;
	assign MC_E_in4_valid = store_0_out1_valid;
	assign store_0_out1_ready = MC_E_in4_ready;
	assign MC_E_in3_data = store_0_out2_data;
	assign MC_E_in3_valid = store_0_out2_valid;
	assign store_0_out2_ready = MC_E_in3_ready;

	assign cst_9_clk = clk;
	assign cst_9_rst = rst;
	assign add_31_in2_data = cst_9_out1_data;
	assign add_31_in2_valid = cst_9_out1_valid;
	assign cst_9_out1_ready = add_31_in2_ready;

	assign add_31_clk = clk;
	assign add_31_rst = rst;
	assign fork_4_in1_data = add_31_out1_data;
	assign fork_4_in1_valid = add_31_out1_valid;
	assign add_31_out1_ready = fork_4_in1_ready;

	assign cst_10_clk = clk;
	assign cst_10_rst = rst;
	assign icmp_32_in2_data = cst_10_out1_data;
	assign icmp_32_in2_valid = cst_10_out1_valid;
	assign cst_10_out1_ready = icmp_32_in2_ready;

	assign icmp_32_clk = clk;
	assign icmp_32_rst = rst;
	assign fork_37_in1_data = icmp_32_out1_data;
	assign fork_37_in1_valid = icmp_32_out1_valid;
	assign icmp_32_out1_ready = fork_37_in1_ready;

	assign phi_n5_clk = clk;
	assign phi_n5_rst = rst;
	assign fork_21_in1_data = phi_n5_out1_data;
	assign fork_21_in1_valid = phi_n5_out1_valid;
	assign phi_n5_out1_ready = fork_21_in1_ready;

	assign phi_n6_clk = clk;
	assign phi_n6_rst = rst;
	assign fork_22_in1_data = phi_n6_out1_data;
	assign fork_22_in1_valid = phi_n6_out1_valid;
	assign phi_n6_out1_ready = fork_22_in1_ready;

	assign phi_n7_clk = clk;
	assign phi_n7_rst = rst;
	assign store_0_in1_data = phi_n7_out1_data;
	assign store_0_in1_valid = phi_n7_out1_valid;
	assign phi_n7_out1_ready = store_0_in1_ready;

	assign fork_4_clk = clk;
	assign fork_4_rst = rst;
	assign icmp_32_in1_data = fork_4_out1_data;
	assign icmp_32_in1_valid = fork_4_out1_valid;
	assign fork_4_out1_ready = icmp_32_in1_ready;
	assign branch_11_in1_data = fork_4_out2_data;
	assign branch_11_in1_valid = fork_4_out2_valid;
	assign fork_4_out2_ready = branch_11_in1_ready;

	assign fork_21_clk = clk;
	assign fork_21_rst = rst;
	assign shl_27_in1_data = fork_21_out1_data;
	assign shl_27_in1_valid = fork_21_out1_valid;
	assign fork_21_out1_ready = shl_27_in1_ready;
	assign branch_12_in1_data = fork_21_out2_data;
	assign branch_12_in1_valid = fork_21_out2_valid;
	assign fork_21_out2_ready = branch_12_in1_ready;

	assign fork_22_clk = clk;
	assign fork_22_rst = rst;
	assign add_28_in2_data = fork_22_out1_data;
	assign add_28_in2_valid = fork_22_out1_valid;
	assign fork_22_out1_ready = add_28_in2_ready;
	assign add_31_in1_data = fork_22_out2_data;
	assign add_31_in1_valid = fork_22_out2_valid;
	assign fork_22_out2_ready = add_31_in1_ready;

	assign branch_11_clk = clk;
	assign branch_11_rst = rst;
	assign Buffer_105_in1_data = branch_11_out1_data;
	assign Buffer_105_in1_valid = branch_11_out1_valid;
	assign branch_11_out1_ready = Buffer_105_in1_ready;
	assign sink_8_in1_data = branch_11_out2_data;
	assign sink_8_in1_valid = branch_11_out2_valid;
	assign branch_11_out2_ready = sink_8_in1_ready;

	assign branch_12_clk = clk;
	assign branch_12_rst = rst;
	assign Buffer_106_in1_data = branch_12_out1_data;
	assign Buffer_106_in1_valid = branch_12_out1_valid;
	assign branch_12_out1_ready = Buffer_106_in1_ready;
	assign phi_n3_in1_data = branch_12_out2_data;
	assign phi_n3_in1_valid = branch_12_out2_valid;
	assign branch_12_out2_ready = phi_n3_in1_ready;

	assign fork_37_clk = clk;
	assign fork_37_rst = rst;
	assign branch_12_in2_data = fork_37_out1_data;
	assign branch_12_in2_valid = fork_37_out1_valid;
	assign fork_37_out1_ready = branch_12_in2_ready;
	assign branch_11_in2_data = fork_37_out2_data;
	assign branch_11_in2_valid = fork_37_out2_valid;
	assign fork_37_out2_ready = branch_11_in2_ready;
	assign branchC_46_in2_data = fork_37_out3_data;
	assign branchC_46_in2_valid = fork_37_out3_valid;
	assign fork_37_out3_ready = branchC_46_in2_ready;

	assign cst_39_clk = clk;
	assign cst_39_rst = rst;
	assign MC_E_in1_data = cst_39_out1_data;
	assign MC_E_in1_valid = cst_39_out1_valid;
	assign cst_39_out1_ready = MC_E_in1_ready;

	assign phiC_24_clk = clk;
	assign phiC_24_rst = rst;
	assign forkC_57_in1_data = phiC_24_out1_data;
	assign forkC_57_in1_valid = phiC_24_out1_valid;
	assign phiC_24_out1_ready = forkC_57_in1_ready;

	assign forkC_57_clk = clk;
	assign forkC_57_rst = rst;
	assign cst_39_in1_data = forkC_57_out1_data;
	assign cst_39_in1_valid = forkC_57_out1_valid;
	assign forkC_57_out1_ready = cst_39_in1_ready;
	assign branchC_46_in1_data = forkC_57_out2_data;
	assign branchC_46_in1_valid = forkC_57_out2_valid;
	assign forkC_57_out2_ready = branchC_46_in1_ready;

	assign branchC_46_clk = clk;
	assign branchC_46_rst = rst;
	assign Buffer_107_in1_data = branchC_46_out1_data;
	assign Buffer_107_in1_valid = branchC_46_out1_valid;
	assign branchC_46_out1_ready = Buffer_107_in1_ready;
	assign phiC_25_in1_data = branchC_46_out2_data;
	assign phiC_25_in1_valid = branchC_46_out2_valid;
	assign branchC_46_out2_ready = phiC_25_in1_ready;

	assign source_5_clk = clk;
	assign source_5_rst = rst;
	assign cst_8_in1_data = source_5_out1_data;
	assign cst_8_in1_valid = source_5_out1_valid;
	assign source_5_out1_ready = cst_8_in1_ready;

	assign source_6_clk = clk;
	assign source_6_rst = rst;
	assign cst_9_in1_data = source_6_out1_data;
	assign cst_9_in1_valid = source_6_out1_valid;
	assign source_6_out1_ready = cst_9_in1_ready;

	assign source_7_clk = clk;
	assign source_7_rst = rst;
	assign cst_10_in1_data = source_7_out1_data;
	assign cst_10_in1_valid = source_7_out1_valid;
	assign source_7_out1_ready = cst_10_in1_ready;

	assign brCst_block1_clk = clk;
	assign brCst_block1_rst = rst;
	assign fork_53_in1_data = brCst_block1_out1_data;
	assign fork_53_in1_valid = brCst_block1_out1_valid;
	assign brCst_block1_out1_ready = fork_53_in1_ready;

	assign cst_0_clk = clk;
	assign cst_0_rst = rst;
	assign branch_0_in1_data = cst_0_out1_data;
	assign branch_0_in1_valid = cst_0_out1_valid;
	assign cst_0_out1_ready = branch_0_in1_ready;

	assign branch_0_clk = clk;
	assign branch_0_rst = rst;
	assign phi_1_in2_data = branch_0_out1_data;
	assign phi_1_in2_valid = branch_0_out1_valid;
	assign branch_0_out1_ready = phi_1_in2_ready;
	assign sink_0_in1_data = branch_0_out2_data;
	assign sink_0_in1_valid = branch_0_out2_valid;
	assign branch_0_out2_ready = sink_0_in1_ready;

	assign start_0_clk = clk;
	assign start_0_rst = rst;
	assign start_0_in1_data = start_in;
	assign start_0_in1_valid = start_valid;
	assign start_ready = start_0_in1_ready;
	assign forkC_52_in1_data = start_0_out1_data;
	assign forkC_52_in1_valid = start_0_out1_valid;
	assign start_0_out1_ready = forkC_52_in1_ready;

	assign forkC_52_clk = clk;
	assign forkC_52_rst = rst;
	assign cst_0_in1_data = forkC_52_out1_data;
	assign cst_0_in1_valid = forkC_52_out1_valid;
	assign forkC_52_out1_ready = cst_0_in1_ready;
	assign branchC_42_in1_data = forkC_52_out2_data;
	assign branchC_42_in1_valid = forkC_52_out2_valid;
	assign forkC_52_out2_ready = branchC_42_in1_ready;
	assign brCst_block1_in1_data = forkC_52_out3_data;
	assign brCst_block1_in1_valid = forkC_52_out3_valid;
	assign forkC_52_out3_ready = brCst_block1_in1_ready;

	assign branchC_42_clk = clk;
	assign branchC_42_rst = rst;
	assign phiC_21_in1_data = branchC_42_out1_data;
	assign phiC_21_in1_valid = branchC_42_out1_valid;
	assign branchC_42_out1_ready = phiC_21_in1_ready;
	assign sink_30_in1_data = branchC_42_out2_data;
	assign sink_30_in1_valid = branchC_42_out2_valid;
	assign branchC_42_out2_ready = sink_30_in1_ready;

	assign fork_53_clk = clk;
	assign fork_53_rst = rst;
	assign branch_0_in2_data = fork_53_out1_data;
	assign branch_0_in2_valid = fork_53_out1_valid;
	assign fork_53_out1_ready = branch_0_in2_ready;
	assign branchC_42_in2_data = fork_53_out2_data;
	assign branchC_42_in2_valid = fork_53_out2_valid;
	assign fork_53_out2_ready = branchC_42_in2_ready;

	assign phi_77_clk = clk;
	assign phi_77_rst = rst;
	assign fork_12_in1_data = phi_77_out1_data;
	assign fork_12_in1_valid = phi_77_out1_valid;
	assign phi_77_out1_ready = fork_12_in1_ready;

	assign cst_28_clk = clk;
	assign cst_28_rst = rst;
	assign shl_78_in2_data = cst_28_out1_data;
	assign shl_78_in2_valid = cst_28_out1_valid;
	assign cst_28_out1_ready = shl_78_in2_ready;

	assign shl_78_clk = clk;
	assign shl_78_rst = rst;
	assign add_79_in1_data = shl_78_out1_data;
	assign add_79_in1_valid = shl_78_out1_valid;
	assign shl_78_out1_ready = add_79_in1_ready;

	assign add_79_clk = clk;
	assign add_79_rst = rst;
	assign load_82_in2_data = add_79_out1_data;
	assign load_82_in2_valid = add_79_out1_valid;
	assign add_79_out1_ready = load_82_in2_ready;

	assign load_82_clk = clk;
	assign load_82_rst = rst;
	assign branch_31_in1_data = load_82_out1_data;
	assign branch_31_in1_valid = load_82_out1_valid;
	assign load_82_out1_ready = branch_31_in1_ready;
	assign MC_G_in2_data = load_82_out2_data;
	assign MC_G_in2_valid = load_82_out2_valid;
	assign load_82_out2_ready = MC_G_in2_ready;

	assign brCst_block15_clk = clk;
	assign brCst_block15_rst = rst;
	assign fork_47_in1_data = brCst_block15_out1_data;
	assign fork_47_in1_valid = brCst_block15_out1_valid;
	assign brCst_block15_out1_ready = fork_47_in1_ready;

	assign cst_29_clk = clk;
	assign cst_29_rst = rst;
	assign branch_32_in1_data = cst_29_out1_data;
	assign branch_32_in1_valid = cst_29_out1_valid;
	assign cst_29_out1_ready = branch_32_in1_ready;

	assign phi_n15_clk = clk;
	assign phi_n15_rst = rst;
	assign fork_28_in1_data = phi_n15_out1_data;
	assign fork_28_in1_valid = phi_n15_out1_valid;
	assign phi_n15_out1_ready = fork_28_in1_ready;

	assign fork_12_clk = clk;
	assign fork_12_rst = rst;
	assign add_79_in2_data = fork_12_out1_data;
	assign add_79_in2_valid = fork_12_out1_valid;
	assign fork_12_out1_ready = add_79_in2_ready;
	assign branch_33_in1_data = fork_12_out2_data;
	assign branch_33_in1_valid = fork_12_out2_valid;
	assign fork_12_out2_ready = branch_33_in1_ready;

	assign fork_28_clk = clk;
	assign fork_28_rst = rst;
	assign shl_78_in1_data = fork_28_out1_data;
	assign shl_78_in1_valid = fork_28_out1_valid;
	assign fork_28_out1_ready = shl_78_in1_ready;
	assign branch_34_in1_data = fork_28_out2_data;
	assign branch_34_in1_valid = fork_28_out2_valid;
	assign fork_28_out2_ready = branch_34_in1_ready;

	assign branch_31_clk = clk;
	assign branch_31_rst = rst;
	assign phi_84_in2_data = branch_31_out1_data;
	assign phi_84_in2_valid = branch_31_out1_valid;
	assign branch_31_out1_ready = phi_84_in2_ready;
	assign sink_23_in1_data = branch_31_out2_data;
	assign sink_23_in1_valid = branch_31_out2_valid;
	assign branch_31_out2_ready = sink_23_in1_ready;

	assign branch_32_clk = clk;
	assign branch_32_rst = rst;
	assign phi_85_in2_data = branch_32_out1_data;
	assign phi_85_in2_valid = branch_32_out1_valid;
	assign branch_32_out1_ready = phi_85_in2_ready;
	assign sink_24_in1_data = branch_32_out2_data;
	assign sink_24_in1_valid = branch_32_out2_valid;
	assign branch_32_out2_ready = sink_24_in1_ready;

	assign branch_33_clk = clk;
	assign branch_33_rst = rst;
	assign phi_n20_in1_data = branch_33_out1_data;
	assign phi_n20_in1_valid = branch_33_out1_valid;
	assign branch_33_out1_ready = phi_n20_in1_ready;
	assign sink_25_in1_data = branch_33_out2_data;
	assign sink_25_in1_valid = branch_33_out2_valid;
	assign branch_33_out2_ready = sink_25_in1_ready;

	assign branch_34_clk = clk;
	assign branch_34_rst = rst;
	assign phi_n19_in1_data = branch_34_out1_data;
	assign phi_n19_in1_valid = branch_34_out1_valid;
	assign branch_34_out1_ready = phi_n19_in1_ready;
	assign sink_26_in1_data = branch_34_out2_data;
	assign sink_26_in1_valid = branch_34_out2_valid;
	assign branch_34_out2_ready = sink_26_in1_ready;

	assign fork_47_clk = clk;
	assign fork_47_rst = rst;
	assign branch_34_in2_data = fork_47_out1_data;
	assign branch_34_in2_valid = fork_47_out1_valid;
	assign fork_47_out1_ready = branch_34_in2_ready;
	assign branch_33_in2_data = fork_47_out2_data;
	assign branch_33_in2_valid = fork_47_out2_valid;
	assign fork_47_out2_ready = branch_33_in2_ready;
	assign branch_32_in2_data = fork_47_out3_data;
	assign branch_32_in2_valid = fork_47_out3_valid;
	assign fork_47_out3_ready = branch_32_in2_ready;
	assign branch_31_in2_data = fork_47_out4_data;
	assign branch_31_in2_valid = fork_47_out4_valid;
	assign fork_47_out4_ready = branch_31_in2_ready;
	assign branchC_56_in2_data = fork_47_out5_data;
	assign branchC_56_in2_valid = fork_47_out5_valid;
	assign fork_47_out5_ready = branchC_56_in2_ready;

	assign phiC_34_clk = clk;
	assign phiC_34_rst = rst;
	assign forkC_71_in1_data = phiC_34_out1_data;
	assign forkC_71_in1_valid = phiC_34_out1_valid;
	assign phiC_34_out1_ready = forkC_71_in1_ready;
	assign phi_77_in1_data = phiC_34_out2_data;
	assign phi_77_in1_valid = phiC_34_out2_valid;
	assign phiC_34_out2_ready = phi_77_in1_ready;

	assign forkC_71_clk = clk;
	assign forkC_71_rst = rst;
	assign cst_29_in1_data = forkC_71_out1_data;
	assign cst_29_in1_valid = forkC_71_out1_valid;
	assign forkC_71_out1_ready = cst_29_in1_ready;
	assign branchC_56_in1_data = forkC_71_out2_data;
	assign branchC_56_in1_valid = forkC_71_out2_valid;
	assign forkC_71_out2_ready = branchC_56_in1_ready;
	assign brCst_block15_in1_data = forkC_71_out3_data;
	assign brCst_block15_in1_valid = forkC_71_out3_valid;
	assign forkC_71_out3_ready = brCst_block15_in1_ready;

	assign branchC_56_clk = clk;
	assign branchC_56_rst = rst;
	assign phiC_35_in1_data = branchC_56_out1_data;
	assign phiC_35_in1_valid = branchC_56_out1_valid;
	assign branchC_56_out1_ready = phiC_35_in1_ready;
	assign sink_38_in1_data = branchC_56_out2_data;
	assign sink_38_in1_valid = branchC_56_out2_valid;
	assign branchC_56_out2_ready = sink_38_in1_ready;

	assign source_20_clk = clk;
	assign source_20_rst = rst;
	assign cst_28_in1_data = source_20_out1_data;
	assign cst_28_in1_valid = source_20_out1_valid;
	assign source_20_out1_ready = cst_28_in1_ready;

	assign phi_38_clk = clk;
	assign phi_38_rst = rst;
	assign branch_16_in1_data = phi_38_out1_data;
	assign branch_16_in1_valid = phi_38_out1_valid;
	assign phi_38_out1_ready = branch_16_in1_ready;

	assign brCst_block8_clk = clk;
	assign brCst_block8_rst = rst;
	assign fork_40_in1_data = brCst_block8_out1_data;
	assign fork_40_in1_valid = brCst_block8_out1_valid;
	assign brCst_block8_out1_ready = fork_40_in1_ready;

	assign cst_14_clk = clk;
	assign cst_14_rst = rst;
	assign branch_15_in1_data = cst_14_out1_data;
	assign branch_15_in1_valid = cst_14_out1_valid;
	assign cst_14_out1_ready = branch_15_in1_ready;

	assign branch_15_clk = clk;
	assign branch_15_rst = rst;
	assign phi_40_in2_data = branch_15_out1_data;
	assign phi_40_in2_valid = branch_15_out1_valid;
	assign branch_15_out1_ready = phi_40_in2_ready;
	assign sink_11_in1_data = branch_15_out2_data;
	assign sink_11_in1_valid = branch_15_out2_valid;
	assign branch_15_out2_ready = sink_11_in1_ready;

	assign branch_16_clk = clk;
	assign branch_16_rst = rst;
	assign phi_n13_in1_data = branch_16_out1_data;
	assign phi_n13_in1_valid = branch_16_out1_valid;
	assign branch_16_out1_ready = phi_n13_in1_ready;
	assign sink_12_in1_data = branch_16_out2_data;
	assign sink_12_in1_valid = branch_16_out2_valid;
	assign branch_16_out2_ready = sink_12_in1_ready;

	assign fork_40_clk = clk;
	assign fork_40_rst = rst;
	assign branch_16_in2_data = fork_40_out1_data;
	assign branch_16_in2_valid = fork_40_out1_valid;
	assign fork_40_out1_ready = branch_16_in2_ready;
	assign branch_15_in2_data = fork_40_out2_data;
	assign branch_15_in2_valid = fork_40_out2_valid;
	assign fork_40_out2_ready = branch_15_in2_ready;
	assign branchC_49_in2_data = fork_40_out3_data;
	assign branchC_49_in2_valid = fork_40_out3_valid;
	assign fork_40_out3_ready = branchC_49_in2_ready;

	assign phiC_27_clk = clk;
	assign phiC_27_rst = rst;
	assign forkC_62_in1_data = phiC_27_out1_data;
	assign forkC_62_in1_valid = phiC_27_out1_valid;
	assign phiC_27_out1_ready = forkC_62_in1_ready;
	assign phi_38_in1_data = phiC_27_out2_data;
	assign phi_38_in1_valid = phiC_27_out2_valid;
	assign phiC_27_out2_ready = phi_38_in1_ready;

	assign forkC_62_clk = clk;
	assign forkC_62_rst = rst;
	assign cst_14_in1_data = forkC_62_out1_data;
	assign cst_14_in1_valid = forkC_62_out1_valid;
	assign forkC_62_out1_ready = cst_14_in1_ready;
	assign branchC_49_in1_data = forkC_62_out2_data;
	assign branchC_49_in1_valid = forkC_62_out2_valid;
	assign forkC_62_out2_ready = branchC_49_in1_ready;
	assign brCst_block8_in1_data = forkC_62_out3_data;
	assign brCst_block8_in1_valid = forkC_62_out3_valid;
	assign forkC_62_out3_ready = brCst_block8_in1_ready;

	assign branchC_49_clk = clk;
	assign branchC_49_rst = rst;
	assign phiC_28_in1_data = branchC_49_out1_data;
	assign phiC_28_in1_valid = branchC_49_out1_valid;
	assign branchC_49_out1_ready = phiC_28_in1_ready;
	assign sink_34_in1_data = branchC_49_out2_data;
	assign sink_34_in1_valid = branchC_49_out2_valid;
	assign branchC_49_out2_ready = sink_34_in1_ready;

	assign cst_11_clk = clk;
	assign cst_11_rst = rst;
	assign add_34_in2_data = cst_11_out1_data;
	assign add_34_in2_valid = cst_11_out1_valid;
	assign cst_11_out1_ready = add_34_in2_ready;

	assign add_34_clk = clk;
	assign add_34_rst = rst;
	assign fork_5_in1_data = add_34_out1_data;
	assign fork_5_in1_valid = add_34_out1_valid;
	assign add_34_out1_ready = fork_5_in1_ready;

	assign cst_12_clk = clk;
	assign cst_12_rst = rst;
	assign icmp_35_in2_data = cst_12_out1_data;
	assign icmp_35_in2_valid = cst_12_out1_valid;
	assign cst_12_out1_ready = icmp_35_in2_ready;

	assign icmp_35_clk = clk;
	assign icmp_35_rst = rst;
	assign fork_59_in1_data = icmp_35_out1_data;
	assign fork_59_in1_valid = icmp_35_out1_valid;
	assign icmp_35_out1_ready = fork_59_in1_ready;

	assign phi_n3_clk = clk;
	assign phi_n3_rst = rst;
	assign add_34_in1_data = phi_n3_out1_data;
	assign add_34_in1_valid = phi_n3_out1_valid;
	assign phi_n3_out1_ready = add_34_in1_ready;

	assign fork_5_clk = clk;
	assign fork_5_rst = rst;
	assign icmp_35_in1_data = fork_5_out1_data;
	assign icmp_35_in1_valid = fork_5_out1_valid;
	assign fork_5_out1_ready = icmp_35_in1_ready;
	assign branch_13_in1_data = fork_5_out2_data;
	assign branch_13_in1_valid = fork_5_out2_valid;
	assign fork_5_out2_ready = branch_13_in1_ready;

	assign branch_13_clk = clk;
	assign branch_13_rst = rst;
	assign Buffer_108_in1_data = branch_13_out1_data;
	assign Buffer_108_in1_valid = branch_13_out1_valid;
	assign branch_13_out1_ready = Buffer_108_in1_ready;
	assign sink_9_in1_data = branch_13_out2_data;
	assign sink_9_in1_valid = branch_13_out2_valid;
	assign branch_13_out2_ready = sink_9_in1_ready;

	assign phiC_25_clk = clk;
	assign phiC_25_rst = rst;
	assign branchC_47_in1_data = phiC_25_out1_data;
	assign branchC_47_in1_valid = phiC_25_out1_valid;
	assign phiC_25_out1_ready = branchC_47_in1_ready;

	assign branchC_47_clk = clk;
	assign branchC_47_rst = rst;
	assign Buffer_109_in1_data = branchC_47_out1_data;
	assign Buffer_109_in1_valid = branchC_47_out1_valid;
	assign branchC_47_out1_ready = Buffer_109_in1_ready;
	assign phiC_26_in1_data = branchC_47_out2_data;
	assign phiC_26_in1_valid = branchC_47_out2_valid;
	assign branchC_47_out2_ready = phiC_26_in1_ready;

	assign fork_59_clk = clk;
	assign fork_59_rst = rst;
	assign branch_13_in2_data = fork_59_out1_data;
	assign branch_13_in2_valid = fork_59_out1_valid;
	assign fork_59_out1_ready = branch_13_in2_ready;
	assign branchC_47_in2_data = fork_59_out2_data;
	assign branchC_47_in2_valid = fork_59_out2_valid;
	assign fork_59_out2_ready = branchC_47_in2_ready;

	assign source_8_clk = clk;
	assign source_8_rst = rst;
	assign cst_11_in1_data = source_8_out1_data;
	assign cst_11_in1_valid = source_8_out1_valid;
	assign source_8_out1_ready = cst_11_in1_ready;

	assign source_9_clk = clk;
	assign source_9_rst = rst;
	assign cst_12_in1_data = source_9_out1_data;
	assign cst_12_in1_valid = source_9_out1_valid;
	assign source_9_out1_ready = cst_12_in1_ready;

	assign cst_34_clk = clk;
	assign cst_34_rst = rst;
	assign shl_101_in2_data = cst_34_out1_data;
	assign shl_101_in2_valid = cst_34_out1_valid;
	assign cst_34_out1_ready = shl_101_in2_ready;

	assign shl_101_clk = clk;
	assign shl_101_rst = rst;
	assign add_102_in1_data = shl_101_out1_data;
	assign add_102_in1_valid = shl_101_out1_valid;
	assign shl_101_out1_ready = add_102_in1_ready;

	assign add_102_clk = clk;
	assign add_102_rst = rst;
	assign store_2_in2_data = add_102_out1_data;
	assign store_2_in2_valid = add_102_out1_valid;
	assign add_102_out1_ready = store_2_in2_ready;

	assign store_2_clk = clk;
	assign store_2_rst = rst;
	assign MC_G_in4_data = store_2_out1_data;
	assign MC_G_in4_valid = store_2_out1_valid;
	assign store_2_out1_ready = MC_G_in4_ready;
	assign MC_G_in3_data = store_2_out2_data;
	assign MC_G_in3_valid = store_2_out2_valid;
	assign store_2_out2_ready = MC_G_in3_ready;

	assign cst_35_clk = clk;
	assign cst_35_rst = rst;
	assign add_105_in2_data = cst_35_out1_data;
	assign add_105_in2_valid = cst_35_out1_valid;
	assign cst_35_out1_ready = add_105_in2_ready;

	assign add_105_clk = clk;
	assign add_105_rst = rst;
	assign fork_16_in1_data = add_105_out1_data;
	assign fork_16_in1_valid = add_105_out1_valid;
	assign add_105_out1_ready = fork_16_in1_ready;

	assign cst_36_clk = clk;
	assign cst_36_rst = rst;
	assign icmp_106_in2_data = cst_36_out1_data;
	assign icmp_106_in2_valid = cst_36_out1_valid;
	assign cst_36_out1_ready = icmp_106_in2_ready;

	assign icmp_106_clk = clk;
	assign icmp_106_rst = rst;
	assign fork_49_in1_data = icmp_106_out1_data;
	assign fork_49_in1_valid = icmp_106_out1_valid;
	assign icmp_106_out1_ready = fork_49_in1_ready;

	assign phi_n16_clk = clk;
	assign phi_n16_rst = rst;
	assign fork_29_in1_data = phi_n16_out1_data;
	assign fork_29_in1_valid = phi_n16_out1_valid;
	assign phi_n16_out1_ready = fork_29_in1_ready;

	assign phi_n17_clk = clk;
	assign phi_n17_rst = rst;
	assign fork_30_in1_data = phi_n17_out1_data;
	assign fork_30_in1_valid = phi_n17_out1_valid;
	assign phi_n17_out1_ready = fork_30_in1_ready;

	assign phi_n18_clk = clk;
	assign phi_n18_rst = rst;
	assign store_2_in1_data = phi_n18_out1_data;
	assign store_2_in1_valid = phi_n18_out1_valid;
	assign phi_n18_out1_ready = store_2_in1_ready;

	assign fork_16_clk = clk;
	assign fork_16_rst = rst;
	assign icmp_106_in1_data = fork_16_out1_data;
	assign icmp_106_in1_valid = fork_16_out1_valid;
	assign fork_16_out1_ready = icmp_106_in1_ready;
	assign branch_39_in1_data = fork_16_out2_data;
	assign branch_39_in1_valid = fork_16_out2_valid;
	assign fork_16_out2_ready = branch_39_in1_ready;

	assign fork_29_clk = clk;
	assign fork_29_rst = rst;
	assign shl_101_in1_data = fork_29_out1_data;
	assign shl_101_in1_valid = fork_29_out1_valid;
	assign fork_29_out1_ready = shl_101_in1_ready;
	assign branch_40_in1_data = fork_29_out2_data;
	assign branch_40_in1_valid = fork_29_out2_valid;
	assign fork_29_out2_ready = branch_40_in1_ready;

	assign fork_30_clk = clk;
	assign fork_30_rst = rst;
	assign add_102_in2_data = fork_30_out1_data;
	assign add_102_in2_valid = fork_30_out1_valid;
	assign fork_30_out1_ready = add_102_in2_ready;
	assign add_105_in1_data = fork_30_out2_data;
	assign add_105_in1_valid = fork_30_out2_valid;
	assign fork_30_out2_ready = add_105_in1_ready;

	assign branch_39_clk = clk;
	assign branch_39_rst = rst;
	assign Buffer_125_in1_data = branch_39_out1_data;
	assign Buffer_125_in1_valid = branch_39_out1_valid;
	assign branch_39_out1_ready = Buffer_125_in1_ready;
	assign sink_28_in1_data = branch_39_out2_data;
	assign sink_28_in1_valid = branch_39_out2_valid;
	assign branch_39_out2_ready = sink_28_in1_ready;

	assign branch_40_clk = clk;
	assign branch_40_rst = rst;
	assign Buffer_126_in1_data = branch_40_out1_data;
	assign Buffer_126_in1_valid = branch_40_out1_valid;
	assign branch_40_out1_ready = Buffer_126_in1_ready;
	assign phi_n14_in1_data = branch_40_out2_data;
	assign phi_n14_in1_valid = branch_40_out2_valid;
	assign branch_40_out2_ready = phi_n14_in1_ready;

	assign fork_49_clk = clk;
	assign fork_49_rst = rst;
	assign branch_40_in2_data = fork_49_out1_data;
	assign branch_40_in2_valid = fork_49_out1_valid;
	assign fork_49_out1_ready = branch_40_in2_ready;
	assign branch_39_in2_data = fork_49_out2_data;
	assign branch_39_in2_valid = fork_49_out2_valid;
	assign fork_49_out2_ready = branch_39_in2_ready;
	assign branchC_58_in2_data = fork_49_out3_data;
	assign branchC_58_in2_valid = fork_49_out3_valid;
	assign fork_49_out3_ready = branchC_58_in2_ready;

	assign cst_41_clk = clk;
	assign cst_41_rst = rst;
	assign MC_G_in1_data = cst_41_out1_data;
	assign MC_G_in1_valid = cst_41_out1_valid;
	assign cst_41_out1_ready = MC_G_in1_ready;

	assign phiC_36_clk = clk;
	assign phiC_36_rst = rst;
	assign forkC_73_in1_data = phiC_36_out1_data;
	assign forkC_73_in1_valid = phiC_36_out1_valid;
	assign phiC_36_out1_ready = forkC_73_in1_ready;

	assign forkC_73_clk = clk;
	assign forkC_73_rst = rst;
	assign cst_41_in1_data = forkC_73_out1_data;
	assign cst_41_in1_valid = forkC_73_out1_valid;
	assign forkC_73_out1_ready = cst_41_in1_ready;
	assign branchC_58_in1_data = forkC_73_out2_data;
	assign branchC_58_in1_valid = forkC_73_out2_valid;
	assign forkC_73_out2_ready = branchC_58_in1_ready;

	assign branchC_58_clk = clk;
	assign branchC_58_rst = rst;
	assign Buffer_127_in1_data = branchC_58_out1_data;
	assign Buffer_127_in1_valid = branchC_58_out1_valid;
	assign branchC_58_out1_ready = Buffer_127_in1_ready;
	assign phiC_37_in1_data = branchC_58_out2_data;
	assign phiC_37_in1_valid = branchC_58_out2_valid;
	assign branchC_58_out2_ready = phiC_37_in1_ready;

	assign source_25_clk = clk;
	assign source_25_rst = rst;
	assign cst_34_in1_data = source_25_out1_data;
	assign cst_34_in1_valid = source_25_out1_valid;
	assign source_25_out1_ready = cst_34_in1_ready;

	assign source_26_clk = clk;
	assign source_26_rst = rst;
	assign cst_35_in1_data = source_26_out1_data;
	assign cst_35_in1_valid = source_26_out1_valid;
	assign source_26_out1_ready = cst_35_in1_ready;

	assign source_27_clk = clk;
	assign source_27_rst = rst;
	assign cst_36_in1_data = source_27_out1_data;
	assign cst_36_in1_valid = source_27_out1_valid;
	assign source_27_out1_ready = cst_36_in1_ready;

	assign cst_21_clk = clk;
	assign cst_21_rst = rst;
	assign shl_64_in2_data = cst_21_out1_data;
	assign shl_64_in2_valid = cst_21_out1_valid;
	assign cst_21_out1_ready = shl_64_in2_ready;

	assign shl_64_clk = clk;
	assign shl_64_rst = rst;
	assign add_65_in1_data = shl_64_out1_data;
	assign add_65_in1_valid = shl_64_out1_valid;
	assign shl_64_out1_ready = add_65_in1_ready;

	assign add_65_clk = clk;
	assign add_65_rst = rst;
	assign store_1_in2_data = add_65_out1_data;
	assign store_1_in2_valid = add_65_out1_valid;
	assign add_65_out1_ready = store_1_in2_ready;

	assign store_1_clk = clk;
	assign store_1_rst = rst;
	assign MC_F_in4_data = store_1_out1_data;
	assign MC_F_in4_valid = store_1_out1_valid;
	assign store_1_out1_ready = MC_F_in4_ready;
	assign MC_F_in3_data = store_1_out2_data;
	assign MC_F_in3_valid = store_1_out2_valid;
	assign store_1_out2_ready = MC_F_in3_ready;

	assign cst_22_clk = clk;
	assign cst_22_rst = rst;
	assign add_68_in2_data = cst_22_out1_data;
	assign add_68_in2_valid = cst_22_out1_valid;
	assign cst_22_out1_ready = add_68_in2_ready;

	assign add_68_clk = clk;
	assign add_68_rst = rst;
	assign fork_10_in1_data = add_68_out1_data;
	assign fork_10_in1_valid = add_68_out1_valid;
	assign add_68_out1_ready = fork_10_in1_ready;

	assign cst_23_clk = clk;
	assign cst_23_rst = rst;
	assign icmp_69_in2_data = cst_23_out1_data;
	assign icmp_69_in2_valid = cst_23_out1_valid;
	assign cst_23_out1_ready = icmp_69_in2_ready;

	assign icmp_69_clk = clk;
	assign icmp_69_rst = rst;
	assign fork_43_in1_data = icmp_69_out1_data;
	assign fork_43_in1_valid = icmp_69_out1_valid;
	assign icmp_69_out1_ready = fork_43_in1_ready;

	assign phi_n0_clk = clk;
	assign phi_n0_rst = rst;
	assign fork_18_in1_data = phi_n0_out1_data;
	assign fork_18_in1_valid = phi_n0_out1_valid;
	assign phi_n0_out1_ready = fork_18_in1_ready;

	assign phi_n1_clk = clk;
	assign phi_n1_rst = rst;
	assign fork_19_in1_data = phi_n1_out1_data;
	assign fork_19_in1_valid = phi_n1_out1_valid;
	assign phi_n1_out1_ready = fork_19_in1_ready;

	assign phi_n2_clk = clk;
	assign phi_n2_rst = rst;
	assign store_1_in1_data = phi_n2_out1_data;
	assign store_1_in1_valid = phi_n2_out1_valid;
	assign phi_n2_out1_ready = store_1_in1_ready;

	assign fork_10_clk = clk;
	assign fork_10_rst = rst;
	assign icmp_69_in1_data = fork_10_out1_data;
	assign icmp_69_in1_valid = fork_10_out1_valid;
	assign fork_10_out1_ready = icmp_69_in1_ready;
	assign branch_25_in1_data = fork_10_out2_data;
	assign branch_25_in1_valid = fork_10_out2_valid;
	assign fork_10_out2_ready = branch_25_in1_ready;

	assign fork_18_clk = clk;
	assign fork_18_rst = rst;
	assign shl_64_in1_data = fork_18_out1_data;
	assign shl_64_in1_valid = fork_18_out1_valid;
	assign fork_18_out1_ready = shl_64_in1_ready;
	assign branch_26_in1_data = fork_18_out2_data;
	assign branch_26_in1_valid = fork_18_out2_valid;
	assign fork_18_out2_ready = branch_26_in1_ready;

	assign fork_19_clk = clk;
	assign fork_19_rst = rst;
	assign add_65_in2_data = fork_19_out1_data;
	assign add_65_in2_valid = fork_19_out1_valid;
	assign fork_19_out1_ready = add_65_in2_ready;
	assign add_68_in1_data = fork_19_out2_data;
	assign add_68_in1_valid = fork_19_out2_valid;
	assign fork_19_out2_ready = add_68_in1_ready;

	assign branch_25_clk = clk;
	assign branch_25_rst = rst;
	assign Buffer_115_in1_data = branch_25_out1_data;
	assign Buffer_115_in1_valid = branch_25_out1_valid;
	assign branch_25_out1_ready = Buffer_115_in1_ready;
	assign sink_18_in1_data = branch_25_out2_data;
	assign sink_18_in1_valid = branch_25_out2_valid;
	assign branch_25_out2_ready = sink_18_in1_ready;

	assign branch_26_clk = clk;
	assign branch_26_rst = rst;
	assign Buffer_116_in1_data = branch_26_out1_data;
	assign Buffer_116_in1_valid = branch_26_out1_valid;
	assign branch_26_out1_ready = Buffer_116_in1_ready;
	assign phi_n12_in1_data = branch_26_out2_data;
	assign phi_n12_in1_valid = branch_26_out2_valid;
	assign branch_26_out2_ready = phi_n12_in1_ready;

	assign fork_43_clk = clk;
	assign fork_43_rst = rst;
	assign branch_26_in2_data = fork_43_out1_data;
	assign branch_26_in2_valid = fork_43_out1_valid;
	assign fork_43_out1_ready = branch_26_in2_ready;
	assign branch_25_in2_data = fork_43_out2_data;
	assign branch_25_in2_valid = fork_43_out2_valid;
	assign fork_43_out2_ready = branch_25_in2_ready;
	assign branchC_52_in2_data = fork_43_out3_data;
	assign branchC_52_in2_valid = fork_43_out3_valid;
	assign fork_43_out3_ready = branchC_52_in2_ready;

	assign cst_40_clk = clk;
	assign cst_40_rst = rst;
	assign MC_F_in1_data = cst_40_out1_data;
	assign MC_F_in1_valid = cst_40_out1_valid;
	assign cst_40_out1_ready = MC_F_in1_ready;

	assign phiC_30_clk = clk;
	assign phiC_30_rst = rst;
	assign forkC_65_in1_data = phiC_30_out1_data;
	assign forkC_65_in1_valid = phiC_30_out1_valid;
	assign phiC_30_out1_ready = forkC_65_in1_ready;

	assign forkC_65_clk = clk;
	assign forkC_65_rst = rst;
	assign cst_40_in1_data = forkC_65_out1_data;
	assign cst_40_in1_valid = forkC_65_out1_valid;
	assign forkC_65_out1_ready = cst_40_in1_ready;
	assign branchC_52_in1_data = forkC_65_out2_data;
	assign branchC_52_in1_valid = forkC_65_out2_valid;
	assign forkC_65_out2_ready = branchC_52_in1_ready;

	assign branchC_52_clk = clk;
	assign branchC_52_rst = rst;
	assign Buffer_117_in1_data = branchC_52_out1_data;
	assign Buffer_117_in1_valid = branchC_52_out1_valid;
	assign branchC_52_out1_ready = Buffer_117_in1_ready;
	assign phiC_31_in1_data = branchC_52_out2_data;
	assign phiC_31_in1_valid = branchC_52_out2_valid;
	assign branchC_52_out2_ready = phiC_31_in1_ready;

	assign source_15_clk = clk;
	assign source_15_rst = rst;
	assign cst_21_in1_data = source_15_out1_data;
	assign cst_21_in1_valid = source_15_out1_valid;
	assign source_15_out1_ready = cst_21_in1_ready;

	assign source_16_clk = clk;
	assign source_16_rst = rst;
	assign cst_22_in1_data = source_16_out1_data;
	assign cst_22_in1_valid = source_16_out1_valid;
	assign source_16_out1_ready = cst_22_in1_ready;

	assign source_17_clk = clk;
	assign source_17_rst = rst;
	assign cst_23_in1_data = source_17_out1_data;
	assign cst_23_in1_valid = source_17_out1_valid;
	assign source_17_out1_ready = cst_23_in1_ready;

	assign phi_40_clk = clk;
	assign phi_40_rst = rst;
	assign fork_6_in1_data = phi_40_out1_data;
	assign fork_6_in1_valid = phi_40_out1_valid;
	assign phi_40_out1_ready = fork_6_in1_ready;

	assign cst_15_clk = clk;
	assign cst_15_rst = rst;
	assign shl_41_in2_data = cst_15_out1_data;
	assign shl_41_in2_valid = cst_15_out1_valid;
	assign cst_15_out1_ready = shl_41_in2_ready;

	assign shl_41_clk = clk;
	assign shl_41_rst = rst;
	assign add_42_in1_data = shl_41_out1_data;
	assign add_42_in1_valid = shl_41_out1_valid;
	assign shl_41_out1_ready = add_42_in1_ready;

	assign add_42_clk = clk;
	assign add_42_rst = rst;
	assign load_45_in2_data = add_42_out1_data;
	assign load_45_in2_valid = add_42_out1_valid;
	assign add_42_out1_ready = load_45_in2_ready;

	assign load_45_clk = clk;
	assign load_45_rst = rst;
	assign branch_17_in1_data = load_45_out1_data;
	assign branch_17_in1_valid = load_45_out1_valid;
	assign load_45_out1_ready = branch_17_in1_ready;
	assign MC_F_in2_data = load_45_out2_data;
	assign MC_F_in2_valid = load_45_out2_valid;
	assign load_45_out2_ready = MC_F_in2_ready;

	assign brCst_block9_clk = clk;
	assign brCst_block9_rst = rst;
	assign fork_41_in1_data = brCst_block9_out1_data;
	assign fork_41_in1_valid = brCst_block9_out1_valid;
	assign brCst_block9_out1_ready = fork_41_in1_ready;

	assign cst_16_clk = clk;
	assign cst_16_rst = rst;
	assign branch_18_in1_data = cst_16_out1_data;
	assign branch_18_in1_valid = cst_16_out1_valid;
	assign cst_16_out1_ready = branch_18_in1_ready;

	assign phi_n13_clk = clk;
	assign phi_n13_rst = rst;
	assign fork_27_in1_data = phi_n13_out1_data;
	assign fork_27_in1_valid = phi_n13_out1_valid;
	assign phi_n13_out1_ready = fork_27_in1_ready;

	assign fork_6_clk = clk;
	assign fork_6_rst = rst;
	assign add_42_in2_data = fork_6_out1_data;
	assign add_42_in2_valid = fork_6_out1_valid;
	assign fork_6_out1_ready = add_42_in2_ready;
	assign branch_19_in1_data = fork_6_out2_data;
	assign branch_19_in1_valid = fork_6_out2_valid;
	assign fork_6_out2_ready = branch_19_in1_ready;

	assign fork_27_clk = clk;
	assign fork_27_rst = rst;
	assign shl_41_in1_data = fork_27_out1_data;
	assign shl_41_in1_valid = fork_27_out1_valid;
	assign fork_27_out1_ready = shl_41_in1_ready;
	assign branch_20_in1_data = fork_27_out2_data;
	assign branch_20_in1_valid = fork_27_out2_valid;
	assign fork_27_out2_ready = branch_20_in1_ready;

	assign branch_17_clk = clk;
	assign branch_17_rst = rst;
	assign phi_47_in2_data = branch_17_out1_data;
	assign phi_47_in2_valid = branch_17_out1_valid;
	assign branch_17_out1_ready = phi_47_in2_ready;
	assign sink_13_in1_data = branch_17_out2_data;
	assign sink_13_in1_valid = branch_17_out2_valid;
	assign branch_17_out2_ready = sink_13_in1_ready;

	assign branch_18_clk = clk;
	assign branch_18_rst = rst;
	assign phi_48_in2_data = branch_18_out1_data;
	assign phi_48_in2_valid = branch_18_out1_valid;
	assign branch_18_out1_ready = phi_48_in2_ready;
	assign sink_14_in1_data = branch_18_out2_data;
	assign sink_14_in1_valid = branch_18_out2_valid;
	assign branch_18_out2_ready = sink_14_in1_ready;

	assign branch_19_clk = clk;
	assign branch_19_rst = rst;
	assign phi_n11_in1_data = branch_19_out1_data;
	assign phi_n11_in1_valid = branch_19_out1_valid;
	assign branch_19_out1_ready = phi_n11_in1_ready;
	assign sink_15_in1_data = branch_19_out2_data;
	assign sink_15_in1_valid = branch_19_out2_valid;
	assign branch_19_out2_ready = sink_15_in1_ready;

	assign branch_20_clk = clk;
	assign branch_20_rst = rst;
	assign phi_n10_in1_data = branch_20_out1_data;
	assign phi_n10_in1_valid = branch_20_out1_valid;
	assign branch_20_out1_ready = phi_n10_in1_ready;
	assign sink_16_in1_data = branch_20_out2_data;
	assign sink_16_in1_valid = branch_20_out2_valid;
	assign branch_20_out2_ready = sink_16_in1_ready;

	assign fork_41_clk = clk;
	assign fork_41_rst = rst;
	assign branch_20_in2_data = fork_41_out1_data;
	assign branch_20_in2_valid = fork_41_out1_valid;
	assign fork_41_out1_ready = branch_20_in2_ready;
	assign branch_19_in2_data = fork_41_out2_data;
	assign branch_19_in2_valid = fork_41_out2_valid;
	assign fork_41_out2_ready = branch_19_in2_ready;
	assign branch_18_in2_data = fork_41_out3_data;
	assign branch_18_in2_valid = fork_41_out3_valid;
	assign fork_41_out3_ready = branch_18_in2_ready;
	assign branch_17_in2_data = fork_41_out4_data;
	assign branch_17_in2_valid = fork_41_out4_valid;
	assign fork_41_out4_ready = branch_17_in2_ready;
	assign branchC_50_in2_data = fork_41_out5_data;
	assign branchC_50_in2_valid = fork_41_out5_valid;
	assign fork_41_out5_ready = branchC_50_in2_ready;

	assign phiC_28_clk = clk;
	assign phiC_28_rst = rst;
	assign forkC_63_in1_data = phiC_28_out1_data;
	assign forkC_63_in1_valid = phiC_28_out1_valid;
	assign phiC_28_out1_ready = forkC_63_in1_ready;
	assign phi_40_in1_data = phiC_28_out2_data;
	assign phi_40_in1_valid = phiC_28_out2_valid;
	assign phiC_28_out2_ready = phi_40_in1_ready;

	assign forkC_63_clk = clk;
	assign forkC_63_rst = rst;
	assign cst_16_in1_data = forkC_63_out1_data;
	assign cst_16_in1_valid = forkC_63_out1_valid;
	assign forkC_63_out1_ready = cst_16_in1_ready;
	assign branchC_50_in1_data = forkC_63_out2_data;
	assign branchC_50_in1_valid = forkC_63_out2_valid;
	assign forkC_63_out2_ready = branchC_50_in1_ready;
	assign brCst_block9_in1_data = forkC_63_out3_data;
	assign brCst_block9_in1_valid = forkC_63_out3_valid;
	assign forkC_63_out3_ready = brCst_block9_in1_ready;

	assign branchC_50_clk = clk;
	assign branchC_50_rst = rst;
	assign phiC_29_in1_data = branchC_50_out1_data;
	assign phiC_29_in1_valid = branchC_50_out1_valid;
	assign branchC_50_out1_ready = phiC_29_in1_ready;
	assign sink_35_in1_data = branchC_50_out2_data;
	assign sink_35_in1_valid = branchC_50_out2_valid;
	assign branchC_50_out2_ready = sink_35_in1_ready;

	assign source_10_clk = clk;
	assign source_10_rst = rst;
	assign cst_15_in1_data = source_10_out1_data;
	assign cst_15_in1_valid = source_10_out1_valid;
	assign source_10_out1_ready = cst_15_in1_ready;

	assign brCst_block7_clk = clk;
	assign brCst_block7_rst = rst;
	assign fork_61_in1_data = brCst_block7_out1_data;
	assign fork_61_in1_valid = brCst_block7_out1_valid;
	assign brCst_block7_out1_ready = fork_61_in1_ready;

	assign cst_13_clk = clk;
	assign cst_13_rst = rst;
	assign branch_14_in1_data = cst_13_out1_data;
	assign branch_14_in1_valid = cst_13_out1_valid;
	assign cst_13_out1_ready = branch_14_in1_ready;

	assign branch_14_clk = clk;
	assign branch_14_rst = rst;
	assign phi_38_in2_data = branch_14_out1_data;
	assign phi_38_in2_valid = branch_14_out1_valid;
	assign branch_14_out1_ready = phi_38_in2_ready;
	assign sink_10_in1_data = branch_14_out2_data;
	assign sink_10_in1_valid = branch_14_out2_valid;
	assign branch_14_out2_ready = sink_10_in1_ready;

	assign phiC_26_clk = clk;
	assign phiC_26_rst = rst;
	assign forkC_60_in1_data = phiC_26_out1_data;
	assign forkC_60_in1_valid = phiC_26_out1_valid;
	assign phiC_26_out1_ready = forkC_60_in1_ready;

	assign forkC_60_clk = clk;
	assign forkC_60_rst = rst;
	assign cst_13_in1_data = forkC_60_out1_data;
	assign cst_13_in1_valid = forkC_60_out1_valid;
	assign forkC_60_out1_ready = cst_13_in1_ready;
	assign branchC_48_in1_data = forkC_60_out2_data;
	assign branchC_48_in1_valid = forkC_60_out2_valid;
	assign forkC_60_out2_ready = branchC_48_in1_ready;
	assign brCst_block7_in1_data = forkC_60_out3_data;
	assign brCst_block7_in1_valid = forkC_60_out3_valid;
	assign forkC_60_out3_ready = brCst_block7_in1_ready;

	assign branchC_48_clk = clk;
	assign branchC_48_rst = rst;
	assign phiC_27_in1_data = branchC_48_out1_data;
	assign phiC_27_in1_valid = branchC_48_out1_valid;
	assign branchC_48_out1_ready = phiC_27_in1_ready;
	assign sink_33_in1_data = branchC_48_out2_data;
	assign sink_33_in1_valid = branchC_48_out2_valid;
	assign branchC_48_out2_ready = sink_33_in1_ready;

	assign fork_61_clk = clk;
	assign fork_61_rst = rst;
	assign branch_14_in2_data = fork_61_out1_data;
	assign branch_14_in2_valid = fork_61_out1_valid;
	assign fork_61_out1_ready = branch_14_in2_ready;
	assign branchC_48_in2_data = fork_61_out2_data;
	assign branchC_48_in2_valid = fork_61_out2_valid;
	assign fork_61_out2_ready = branchC_48_in2_ready;

	assign brCst_block13_clk = clk;
	assign brCst_block13_rst = rst;
	assign fork_69_in1_data = brCst_block13_out1_data;
	assign fork_69_in1_valid = brCst_block13_out1_valid;
	assign brCst_block13_out1_ready = fork_69_in1_ready;

	assign cst_26_clk = clk;
	assign cst_26_rst = rst;
	assign branch_28_in1_data = cst_26_out1_data;
	assign branch_28_in1_valid = cst_26_out1_valid;
	assign cst_26_out1_ready = branch_28_in1_ready;

	assign branch_28_clk = clk;
	assign branch_28_rst = rst;
	assign phi_75_in2_data = branch_28_out1_data;
	assign phi_75_in2_valid = branch_28_out1_valid;
	assign branch_28_out1_ready = phi_75_in2_ready;
	assign sink_20_in1_data = branch_28_out2_data;
	assign sink_20_in1_valid = branch_28_out2_valid;
	assign branch_28_out2_ready = sink_20_in1_ready;

	assign phiC_32_clk = clk;
	assign phiC_32_rst = rst;
	assign forkC_68_in1_data = phiC_32_out1_data;
	assign forkC_68_in1_valid = phiC_32_out1_valid;
	assign phiC_32_out1_ready = forkC_68_in1_ready;

	assign forkC_68_clk = clk;
	assign forkC_68_rst = rst;
	assign cst_26_in1_data = forkC_68_out1_data;
	assign cst_26_in1_valid = forkC_68_out1_valid;
	assign forkC_68_out1_ready = cst_26_in1_ready;
	assign branchC_54_in1_data = forkC_68_out2_data;
	assign branchC_54_in1_valid = forkC_68_out2_valid;
	assign forkC_68_out2_ready = branchC_54_in1_ready;
	assign brCst_block13_in1_data = forkC_68_out3_data;
	assign brCst_block13_in1_valid = forkC_68_out3_valid;
	assign forkC_68_out3_ready = brCst_block13_in1_ready;

	assign branchC_54_clk = clk;
	assign branchC_54_rst = rst;
	assign phiC_33_in1_data = branchC_54_out1_data;
	assign phiC_33_in1_valid = branchC_54_out1_valid;
	assign branchC_54_out1_ready = phiC_33_in1_ready;
	assign sink_36_in1_data = branchC_54_out2_data;
	assign sink_36_in1_valid = branchC_54_out2_valid;
	assign branchC_54_out2_ready = sink_36_in1_ready;

	assign fork_69_clk = clk;
	assign fork_69_rst = rst;
	assign branch_28_in2_data = fork_69_out1_data;
	assign branch_28_in2_valid = fork_69_out1_valid;
	assign fork_69_out1_ready = branch_28_in2_ready;
	assign branchC_54_in2_data = fork_69_out2_data;
	assign branchC_54_in2_valid = fork_69_out2_valid;
	assign fork_69_out2_ready = branchC_54_in2_ready;

	assign phi_75_clk = clk;
	assign phi_75_rst = rst;
	assign branch_30_in1_data = phi_75_out1_data;
	assign branch_30_in1_valid = phi_75_out1_valid;
	assign phi_75_out1_ready = branch_30_in1_ready;

	assign brCst_block14_clk = clk;
	assign brCst_block14_rst = rst;
	assign fork_46_in1_data = brCst_block14_out1_data;
	assign fork_46_in1_valid = brCst_block14_out1_valid;
	assign brCst_block14_out1_ready = fork_46_in1_ready;

	assign cst_27_clk = clk;
	assign cst_27_rst = rst;
	assign branch_29_in1_data = cst_27_out1_data;
	assign branch_29_in1_valid = cst_27_out1_valid;
	assign cst_27_out1_ready = branch_29_in1_ready;

	assign branch_29_clk = clk;
	assign branch_29_rst = rst;
	assign phi_77_in2_data = branch_29_out1_data;
	assign phi_77_in2_valid = branch_29_out1_valid;
	assign branch_29_out1_ready = phi_77_in2_ready;
	assign sink_21_in1_data = branch_29_out2_data;
	assign sink_21_in1_valid = branch_29_out2_valid;
	assign branch_29_out2_ready = sink_21_in1_ready;

	assign branch_30_clk = clk;
	assign branch_30_rst = rst;
	assign phi_n15_in1_data = branch_30_out1_data;
	assign phi_n15_in1_valid = branch_30_out1_valid;
	assign branch_30_out1_ready = phi_n15_in1_ready;
	assign sink_22_in1_data = branch_30_out2_data;
	assign sink_22_in1_valid = branch_30_out2_valid;
	assign branch_30_out2_ready = sink_22_in1_ready;

	assign fork_46_clk = clk;
	assign fork_46_rst = rst;
	assign branch_30_in2_data = fork_46_out1_data;
	assign branch_30_in2_valid = fork_46_out1_valid;
	assign fork_46_out1_ready = branch_30_in2_ready;
	assign branch_29_in2_data = fork_46_out2_data;
	assign branch_29_in2_valid = fork_46_out2_valid;
	assign fork_46_out2_ready = branch_29_in2_ready;
	assign branchC_55_in2_data = fork_46_out3_data;
	assign branchC_55_in2_valid = fork_46_out3_valid;
	assign fork_46_out3_ready = branchC_55_in2_ready;

	assign phiC_33_clk = clk;
	assign phiC_33_rst = rst;
	assign forkC_70_in1_data = phiC_33_out1_data;
	assign forkC_70_in1_valid = phiC_33_out1_valid;
	assign phiC_33_out1_ready = forkC_70_in1_ready;
	assign phi_75_in1_data = phiC_33_out2_data;
	assign phi_75_in1_valid = phiC_33_out2_valid;
	assign phiC_33_out2_ready = phi_75_in1_ready;

	assign forkC_70_clk = clk;
	assign forkC_70_rst = rst;
	assign cst_27_in1_data = forkC_70_out1_data;
	assign cst_27_in1_valid = forkC_70_out1_valid;
	assign forkC_70_out1_ready = cst_27_in1_ready;
	assign branchC_55_in1_data = forkC_70_out2_data;
	assign branchC_55_in1_valid = forkC_70_out2_valid;
	assign forkC_70_out2_ready = branchC_55_in1_ready;
	assign brCst_block14_in1_data = forkC_70_out3_data;
	assign brCst_block14_in1_valid = forkC_70_out3_valid;
	assign forkC_70_out3_ready = brCst_block14_in1_ready;

	assign branchC_55_clk = clk;
	assign branchC_55_rst = rst;
	assign phiC_34_in1_data = branchC_55_out1_data;
	assign phiC_34_in1_valid = branchC_55_out1_valid;
	assign branchC_55_out1_ready = phiC_34_in1_ready;
	assign sink_37_in1_data = branchC_55_out2_data;
	assign sink_37_in1_valid = branchC_55_out2_valid;
	assign branchC_55_out2_ready = sink_37_in1_ready;

	assign cst_37_clk = clk;
	assign cst_37_rst = rst;
	assign add_108_in2_data = cst_37_out1_data;
	assign add_108_in2_valid = cst_37_out1_valid;
	assign cst_37_out1_ready = add_108_in2_ready;

	assign add_108_clk = clk;
	assign add_108_rst = rst;
	assign fork_17_in1_data = add_108_out1_data;
	assign fork_17_in1_valid = add_108_out1_valid;
	assign add_108_out1_ready = fork_17_in1_ready;

	assign cst_38_clk = clk;
	assign cst_38_rst = rst;
	assign icmp_109_in2_data = cst_38_out1_data;
	assign icmp_109_in2_valid = cst_38_out1_valid;
	assign cst_38_out1_ready = icmp_109_in2_ready;

	assign icmp_109_clk = clk;
	assign icmp_109_rst = rst;
	assign fork_75_in1_data = icmp_109_out1_data;
	assign fork_75_in1_valid = icmp_109_out1_valid;
	assign icmp_109_out1_ready = fork_75_in1_ready;

	assign phi_n14_clk = clk;
	assign phi_n14_rst = rst;
	assign add_108_in1_data = phi_n14_out1_data;
	assign add_108_in1_valid = phi_n14_out1_valid;
	assign phi_n14_out1_ready = add_108_in1_ready;

	assign fork_17_clk = clk;
	assign fork_17_rst = rst;
	assign icmp_109_in1_data = fork_17_out1_data;
	assign icmp_109_in1_valid = fork_17_out1_valid;
	assign fork_17_out1_ready = icmp_109_in1_ready;
	assign branch_41_in1_data = fork_17_out2_data;
	assign branch_41_in1_valid = fork_17_out2_valid;
	assign fork_17_out2_ready = branch_41_in1_ready;

	assign branch_41_clk = clk;
	assign branch_41_rst = rst;
	assign Buffer_128_in1_data = branch_41_out1_data;
	assign Buffer_128_in1_valid = branch_41_out1_valid;
	assign branch_41_out1_ready = Buffer_128_in1_ready;
	assign sink_29_in1_data = branch_41_out2_data;
	assign sink_29_in1_valid = branch_41_out2_valid;
	assign branch_41_out2_ready = sink_29_in1_ready;

	assign phiC_37_clk = clk;
	assign phiC_37_rst = rst;
	assign branchC_59_in1_data = phiC_37_out1_data;
	assign branchC_59_in1_valid = phiC_37_out1_valid;
	assign phiC_37_out1_ready = branchC_59_in1_ready;

	assign branchC_59_clk = clk;
	assign branchC_59_rst = rst;
	assign Buffer_129_in1_data = branchC_59_out1_data;
	assign Buffer_129_in1_valid = branchC_59_out1_valid;
	assign branchC_59_out1_ready = Buffer_129_in1_ready;
	assign phiC_38_in1_data = branchC_59_out2_data;
	assign phiC_38_in1_valid = branchC_59_out2_valid;
	assign branchC_59_out2_ready = phiC_38_in1_ready;

	assign fork_75_clk = clk;
	assign fork_75_rst = rst;
	assign branch_41_in2_data = fork_75_out1_data;
	assign branch_41_in2_valid = fork_75_out1_valid;
	assign fork_75_out1_ready = branch_41_in2_ready;
	assign branchC_59_in2_data = fork_75_out2_data;
	assign branchC_59_in2_valid = fork_75_out2_valid;
	assign fork_75_out2_ready = branchC_59_in2_ready;

	assign source_28_clk = clk;
	assign source_28_rst = rst;
	assign cst_37_in1_data = source_28_out1_data;
	assign cst_37_in1_valid = source_28_out1_valid;
	assign source_28_out1_ready = cst_37_in1_ready;

	assign source_29_clk = clk;
	assign source_29_rst = rst;
	assign cst_38_in1_data = source_29_out1_data;
	assign cst_38_in1_valid = source_29_out1_valid;
	assign source_29_out1_ready = cst_38_in1_ready;

	assign ret_0_clk = clk;
	assign ret_0_rst = rst;
	assign end_0_in8_data = ret_0_out1_data;
	assign end_0_in8_valid = ret_0_out1_valid;
	assign ret_0_out1_ready = end_0_in8_ready;

	assign end_0_clk = clk;
	assign end_0_rst = rst;
	assign end_out = end_0_out1_data;
	assign end_0_out1_ready = end_ready;
	assign end_valid = end_0_out1_valid;

	assign phiC_38_clk = clk;
	assign phiC_38_rst = rst;
	assign ret_0_in1_data = phiC_38_out1_data;
	assign ret_0_in1_valid = phiC_38_out1_valid;
	assign phiC_38_out1_ready = ret_0_in1_ready;

	assign cst_24_clk = clk;
	assign cst_24_rst = rst;
	assign add_71_in2_data = cst_24_out1_data;
	assign add_71_in2_valid = cst_24_out1_valid;
	assign cst_24_out1_ready = add_71_in2_ready;

	assign add_71_clk = clk;
	assign add_71_rst = rst;
	assign fork_11_in1_data = add_71_out1_data;
	assign fork_11_in1_valid = add_71_out1_valid;
	assign add_71_out1_ready = fork_11_in1_ready;

	assign cst_25_clk = clk;
	assign cst_25_rst = rst;
	assign icmp_72_in2_data = cst_25_out1_data;
	assign icmp_72_in2_valid = cst_25_out1_valid;
	assign cst_25_out1_ready = icmp_72_in2_ready;

	assign icmp_72_clk = clk;
	assign icmp_72_rst = rst;
	assign fork_67_in1_data = icmp_72_out1_data;
	assign fork_67_in1_valid = icmp_72_out1_valid;
	assign icmp_72_out1_ready = fork_67_in1_ready;

	assign phi_n12_clk = clk;
	assign phi_n12_rst = rst;
	assign add_71_in1_data = phi_n12_out1_data;
	assign add_71_in1_valid = phi_n12_out1_valid;
	assign phi_n12_out1_ready = add_71_in1_ready;

	assign fork_11_clk = clk;
	assign fork_11_rst = rst;
	assign icmp_72_in1_data = fork_11_out1_data;
	assign icmp_72_in1_valid = fork_11_out1_valid;
	assign fork_11_out1_ready = icmp_72_in1_ready;
	assign branch_27_in1_data = fork_11_out2_data;
	assign branch_27_in1_valid = fork_11_out2_valid;
	assign fork_11_out2_ready = branch_27_in1_ready;

	assign branch_27_clk = clk;
	assign branch_27_rst = rst;
	assign Buffer_118_in1_data = branch_27_out1_data;
	assign Buffer_118_in1_valid = branch_27_out1_valid;
	assign branch_27_out1_ready = Buffer_118_in1_ready;
	assign sink_19_in1_data = branch_27_out2_data;
	assign sink_19_in1_valid = branch_27_out2_valid;
	assign branch_27_out2_ready = sink_19_in1_ready;

	assign phiC_31_clk = clk;
	assign phiC_31_rst = rst;
	assign branchC_53_in1_data = phiC_31_out1_data;
	assign branchC_53_in1_valid = phiC_31_out1_valid;
	assign phiC_31_out1_ready = branchC_53_in1_ready;

	assign branchC_53_clk = clk;
	assign branchC_53_rst = rst;
	assign Buffer_119_in1_data = branchC_53_out1_data;
	assign Buffer_119_in1_valid = branchC_53_out1_valid;
	assign branchC_53_out1_ready = Buffer_119_in1_ready;
	assign phiC_32_in1_data = branchC_53_out2_data;
	assign phiC_32_in1_valid = branchC_53_out2_valid;
	assign branchC_53_out2_ready = phiC_32_in1_ready;

	assign fork_67_clk = clk;
	assign fork_67_rst = rst;
	assign branch_27_in2_data = fork_67_out1_data;
	assign branch_27_in2_valid = fork_67_out1_valid;
	assign fork_67_out1_ready = branch_27_in2_ready;
	assign branchC_53_in2_data = fork_67_out2_data;
	assign branchC_53_in2_valid = fork_67_out2_valid;
	assign fork_67_out2_ready = branchC_53_in2_ready;

	assign source_18_clk = clk;
	assign source_18_rst = rst;
	assign cst_24_in1_data = source_18_out1_data;
	assign cst_24_in1_valid = source_18_out1_valid;
	assign source_18_out1_ready = cst_24_in1_ready;

	assign source_19_clk = clk;
	assign source_19_rst = rst;
	assign cst_25_in1_data = source_19_out1_data;
	assign cst_25_in1_valid = source_19_out1_valid;
	assign source_19_out1_ready = cst_25_in1_ready;

	assign phi_47_clk = clk;
	assign phi_47_rst = rst;
	assign and_303_in1_data = phi_47_out1_data;
	assign and_303_in1_valid = phi_47_out1_valid;
	assign phi_47_out1_ready = and_303_in1_ready;

	assign phi_48_clk = clk;
	assign phi_48_rst = rst;
	assign fork_7_in1_data = phi_48_out1_data;
	assign fork_7_in1_valid = phi_48_out1_valid;
	assign phi_48_out1_ready = fork_7_in1_ready;

	assign cst_17_clk = clk;
	assign cst_17_rst = rst;
	assign shl_49_in2_data = cst_17_out1_data;
	assign shl_49_in2_valid = cst_17_out1_valid;
	assign cst_17_out1_ready = shl_49_in2_ready;

	assign shl_49_clk = clk;
	assign shl_49_rst = rst;
	assign add_50_in1_data = shl_49_out1_data;
	assign add_50_in1_valid = shl_49_out1_valid;
	assign shl_49_out1_ready = add_50_in1_ready;

	assign add_50_clk = clk;
	assign add_50_rst = rst;
	assign load_53_in2_data = add_50_out1_data;
	assign load_53_in2_valid = add_50_out1_valid;
	assign add_50_out1_ready = load_53_in2_ready;

	assign load_53_clk = clk;
	assign load_53_rst = rst;
	assign and_302_in1_data = load_53_out1_data;
	assign and_302_in1_valid = load_53_out1_valid;
	assign load_53_out1_ready = and_302_in1_ready;
	assign MC_C_in1_data = load_53_out2_data;
	assign MC_C_in1_valid = load_53_out2_valid;
	assign load_53_out2_ready = MC_C_in1_ready;

	assign cst_18_clk = clk;
	assign cst_18_rst = rst;
	assign shl_54_in2_data = cst_18_out1_data;
	assign shl_54_in2_valid = cst_18_out1_valid;
	assign cst_18_out1_ready = shl_54_in2_ready;

	assign shl_54_clk = clk;
	assign shl_54_rst = rst;
	assign add_55_in1_data = shl_54_out1_data;
	assign add_55_in1_valid = shl_54_out1_valid;
	assign shl_54_out1_ready = add_55_in1_ready;

	assign add_55_clk = clk;
	assign add_55_rst = rst;
	assign load_58_in2_data = add_55_out1_data;
	assign load_58_in2_valid = add_55_out1_valid;
	assign add_55_out1_ready = load_58_in2_ready;

	assign load_58_clk = clk;
	assign load_58_rst = rst;
	assign and_302_in2_data = load_58_out1_data;
	assign and_302_in2_valid = load_58_out1_valid;
	assign load_58_out1_ready = and_302_in2_ready;
	assign MC_D_in1_data = load_58_out2_data;
	assign MC_D_in1_valid = load_58_out2_valid;
	assign load_58_out2_ready = MC_D_in1_ready;

	assign cst_19_clk = clk;
	assign cst_19_rst = rst;
	assign add_61_in2_data = cst_19_out1_data;
	assign add_61_in2_valid = cst_19_out1_valid;
	assign cst_19_out1_ready = add_61_in2_ready;

	assign add_61_clk = clk;
	assign add_61_rst = rst;
	assign fork_9_in1_data = add_61_out1_data;
	assign fork_9_in1_valid = add_61_out1_valid;
	assign add_61_out1_ready = fork_9_in1_ready;

	assign cst_20_clk = clk;
	assign cst_20_rst = rst;
	assign icmp_62_in2_data = cst_20_out1_data;
	assign icmp_62_in2_valid = cst_20_out1_valid;
	assign cst_20_out1_ready = icmp_62_in2_ready;

	assign icmp_62_clk = clk;
	assign icmp_62_rst = rst;
	assign fork_42_in1_data = icmp_62_out1_data;
	assign fork_42_in1_valid = icmp_62_out1_valid;
	assign icmp_62_out1_ready = fork_42_in1_ready;

	assign phi_n10_clk = clk;
	assign phi_n10_rst = rst;
	assign fork_25_in1_data = phi_n10_out1_data;
	assign fork_25_in1_valid = phi_n10_out1_valid;
	assign phi_n10_out1_ready = fork_25_in1_ready;

	assign phi_n11_clk = clk;
	assign phi_n11_rst = rst;
	assign fork_26_in1_data = phi_n11_out1_data;
	assign fork_26_in1_valid = phi_n11_out1_valid;
	assign phi_n11_out1_ready = fork_26_in1_ready;

	assign fork_7_clk = clk;
	assign fork_7_rst = rst;
	assign add_50_in2_data = fork_7_out1_data;
	assign add_50_in2_valid = fork_7_out1_valid;
	assign fork_7_out1_ready = add_50_in2_ready;
	assign shl_54_in1_data = fork_7_out2_data;
	assign shl_54_in1_valid = fork_7_out2_valid;
	assign fork_7_out2_ready = shl_54_in1_ready;
	assign add_61_in1_data = fork_7_out3_data;
	assign add_61_in1_valid = fork_7_out3_valid;
	assign fork_7_out3_ready = add_61_in1_ready;

	assign fork_9_clk = clk;
	assign fork_9_rst = rst;
	assign icmp_62_in1_data = fork_9_out1_data;
	assign icmp_62_in1_valid = fork_9_out1_valid;
	assign fork_9_out1_ready = icmp_62_in1_ready;
	assign branch_22_in1_data = fork_9_out2_data;
	assign branch_22_in1_valid = fork_9_out2_valid;
	assign fork_9_out2_ready = branch_22_in1_ready;

	assign fork_25_clk = clk;
	assign fork_25_rst = rst;
	assign shl_49_in1_data = fork_25_out1_data;
	assign shl_49_in1_valid = fork_25_out1_valid;
	assign fork_25_out1_ready = shl_49_in1_ready;
	assign branch_23_in1_data = fork_25_out2_data;
	assign branch_23_in1_valid = fork_25_out2_valid;
	assign fork_25_out2_ready = branch_23_in1_ready;

	assign fork_26_clk = clk;
	assign fork_26_rst = rst;
	assign add_55_in2_data = fork_26_out1_data;
	assign add_55_in2_valid = fork_26_out1_valid;
	assign fork_26_out1_ready = add_55_in2_ready;
	assign branch_24_in1_data = fork_26_out2_data;
	assign branch_24_in1_valid = fork_26_out2_valid;
	assign fork_26_out2_ready = branch_24_in1_ready;

	assign branch_21_clk = clk;
	assign branch_21_rst = rst;
	assign Buffer_110_in1_data = branch_21_out1_data;
	assign Buffer_110_in1_valid = branch_21_out1_valid;
	assign branch_21_out1_ready = Buffer_110_in1_ready;
	assign phi_n2_in1_data = branch_21_out2_data;
	assign phi_n2_in1_valid = branch_21_out2_valid;
	assign branch_21_out2_ready = phi_n2_in1_ready;

	assign branch_22_clk = clk;
	assign branch_22_rst = rst;
	assign Buffer_111_in1_data = branch_22_out1_data;
	assign Buffer_111_in1_valid = branch_22_out1_valid;
	assign branch_22_out1_ready = Buffer_111_in1_ready;
	assign sink_17_in1_data = branch_22_out2_data;
	assign sink_17_in1_valid = branch_22_out2_valid;
	assign branch_22_out2_ready = sink_17_in1_ready;

	assign branch_23_clk = clk;
	assign branch_23_rst = rst;
	assign Buffer_112_in1_data = branch_23_out1_data;
	assign Buffer_112_in1_valid = branch_23_out1_valid;
	assign branch_23_out1_ready = Buffer_112_in1_ready;
	assign phi_n0_in1_data = branch_23_out2_data;
	assign phi_n0_in1_valid = branch_23_out2_valid;
	assign branch_23_out2_ready = phi_n0_in1_ready;

	assign branch_24_clk = clk;
	assign branch_24_rst = rst;
	assign Buffer_113_in1_data = branch_24_out1_data;
	assign Buffer_113_in1_valid = branch_24_out1_valid;
	assign branch_24_out1_ready = Buffer_113_in1_ready;
	assign phi_n1_in1_data = branch_24_out2_data;
	assign phi_n1_in1_valid = branch_24_out2_valid;
	assign branch_24_out2_ready = phi_n1_in1_ready;

	assign fork_42_clk = clk;
	assign fork_42_rst = rst;
	assign branch_24_in2_data = fork_42_out1_data;
	assign branch_24_in2_valid = fork_42_out1_valid;
	assign fork_42_out1_ready = branch_24_in2_ready;
	assign branch_23_in2_data = fork_42_out2_data;
	assign branch_23_in2_valid = fork_42_out2_valid;
	assign fork_42_out2_ready = branch_23_in2_ready;
	assign branch_22_in2_data = fork_42_out3_data;
	assign branch_22_in2_valid = fork_42_out3_valid;
	assign fork_42_out3_ready = branch_22_in2_ready;
	assign branch_21_in2_data = fork_42_out4_data;
	assign branch_21_in2_valid = fork_42_out4_valid;
	assign fork_42_out4_ready = branch_21_in2_ready;
	assign branchC_51_in2_data = fork_42_out5_data;
	assign branchC_51_in2_valid = fork_42_out5_valid;
	assign fork_42_out5_ready = branchC_51_in2_ready;

	assign phiC_29_clk = clk;
	assign phiC_29_rst = rst;
	assign branchC_51_in1_data = phiC_29_out1_data;
	assign branchC_51_in1_valid = phiC_29_out1_valid;
	assign phiC_29_out1_ready = branchC_51_in1_ready;
	assign fork_82_in1_data = phiC_29_out2_data;
	assign fork_82_in1_valid = phiC_29_out2_valid;
	assign phiC_29_out2_ready = fork_82_in1_ready;

	assign branchC_51_clk = clk;
	assign branchC_51_rst = rst;
	assign Buffer_114_in1_data = branchC_51_out1_data;
	assign Buffer_114_in1_valid = branchC_51_out1_valid;
	assign branchC_51_out1_ready = Buffer_114_in1_ready;
	assign phiC_30_in1_data = branchC_51_out2_data;
	assign phiC_30_in1_valid = branchC_51_out2_valid;
	assign branchC_51_out2_ready = phiC_30_in1_ready;

	assign source_11_clk = clk;
	assign source_11_rst = rst;
	assign cst_17_in1_data = source_11_out1_data;
	assign cst_17_in1_valid = source_11_out1_valid;
	assign source_11_out1_ready = cst_17_in1_ready;

	assign source_12_clk = clk;
	assign source_12_rst = rst;
	assign cst_18_in1_data = source_12_out1_data;
	assign cst_18_in1_valid = source_12_out1_valid;
	assign source_12_out1_ready = cst_18_in1_ready;

	assign source_13_clk = clk;
	assign source_13_rst = rst;
	assign cst_19_in1_data = source_13_out1_data;
	assign cst_19_in1_valid = source_13_out1_valid;
	assign source_13_out1_ready = cst_19_in1_ready;

	assign source_14_clk = clk;
	assign source_14_rst = rst;
	assign cst_20_in1_data = source_14_out1_data;
	assign cst_20_in1_valid = source_14_out1_valid;
	assign source_14_out1_ready = cst_20_in1_ready;

	assign fork_82_clk = clk;
	assign fork_82_rst = rst;
	assign phi_47_in1_data = fork_82_out1_data;
	assign phi_47_in1_valid = fork_82_out1_valid;
	assign fork_82_out1_ready = phi_47_in1_ready;
	assign phi_48_in1_data = fork_82_out2_data;
	assign phi_48_in1_valid = fork_82_out2_valid;
	assign fork_82_out2_ready = phi_48_in1_ready;

	assign phi_10_clk = clk;
	assign phi_10_rst = rst;
	assign and_301_in1_data = phi_10_out1_data;
	assign and_301_in1_valid = phi_10_out1_valid;
	assign phi_10_out1_ready = and_301_in1_ready;

	assign phi_11_clk = clk;
	assign phi_11_rst = rst;
	assign fork_1_in1_data = phi_11_out1_data;
	assign fork_1_in1_valid = phi_11_out1_valid;
	assign phi_11_out1_ready = fork_1_in1_ready;

	assign cst_4_clk = clk;
	assign cst_4_rst = rst;
	assign shl_12_in2_data = cst_4_out1_data;
	assign shl_12_in2_valid = cst_4_out1_valid;
	assign cst_4_out1_ready = shl_12_in2_ready;

	assign shl_12_clk = clk;
	assign shl_12_rst = rst;
	assign add_13_in1_data = shl_12_out1_data;
	assign add_13_in1_valid = shl_12_out1_valid;
	assign shl_12_out1_ready = add_13_in1_ready;

	assign add_13_clk = clk;
	assign add_13_rst = rst;
	assign load_16_in2_data = add_13_out1_data;
	assign load_16_in2_valid = add_13_out1_valid;
	assign add_13_out1_ready = load_16_in2_ready;

	assign load_16_clk = clk;
	assign load_16_rst = rst;
	assign and_300_in1_data = load_16_out1_data;
	assign and_300_in1_valid = load_16_out1_valid;
	assign load_16_out1_ready = and_300_in1_ready;
	assign MC_A_in1_data = load_16_out2_data;
	assign MC_A_in1_valid = load_16_out2_valid;
	assign load_16_out2_ready = MC_A_in1_ready;

	assign cst_5_clk = clk;
	assign cst_5_rst = rst;
	assign shl_17_in2_data = cst_5_out1_data;
	assign shl_17_in2_valid = cst_5_out1_valid;
	assign cst_5_out1_ready = shl_17_in2_ready;

	assign shl_17_clk = clk;
	assign shl_17_rst = rst;
	assign add_18_in1_data = shl_17_out1_data;
	assign add_18_in1_valid = shl_17_out1_valid;
	assign shl_17_out1_ready = add_18_in1_ready;

	assign add_18_clk = clk;
	assign add_18_rst = rst;
	assign load_21_in2_data = add_18_out1_data;
	assign load_21_in2_valid = add_18_out1_valid;
	assign add_18_out1_ready = load_21_in2_ready;

	assign load_21_clk = clk;
	assign load_21_rst = rst;
	assign and_300_in2_data = load_21_out1_data;
	assign and_300_in2_valid = load_21_out1_valid;
	assign load_21_out1_ready = and_300_in2_ready;
	assign MC_B_in1_data = load_21_out2_data;
	assign MC_B_in1_valid = load_21_out2_valid;
	assign load_21_out2_ready = MC_B_in1_ready;

	assign cst_6_clk = clk;
	assign cst_6_rst = rst;
	assign add_24_in2_data = cst_6_out1_data;
	assign add_24_in2_valid = cst_6_out1_valid;
	assign cst_6_out1_ready = add_24_in2_ready;

	assign add_24_clk = clk;
	assign add_24_rst = rst;
	assign fork_3_in1_data = add_24_out1_data;
	assign fork_3_in1_valid = add_24_out1_valid;
	assign add_24_out1_ready = fork_3_in1_ready;

	assign cst_7_clk = clk;
	assign cst_7_rst = rst;
	assign icmp_25_in2_data = cst_7_out1_data;
	assign icmp_25_in2_valid = cst_7_out1_valid;
	assign cst_7_out1_ready = icmp_25_in2_ready;

	assign icmp_25_clk = clk;
	assign icmp_25_rst = rst;
	assign fork_36_in1_data = icmp_25_out1_data;
	assign fork_36_in1_valid = icmp_25_out1_valid;
	assign icmp_25_out1_ready = fork_36_in1_ready;

	assign phi_n8_clk = clk;
	assign phi_n8_rst = rst;
	assign fork_23_in1_data = phi_n8_out1_data;
	assign fork_23_in1_valid = phi_n8_out1_valid;
	assign phi_n8_out1_ready = fork_23_in1_ready;

	assign phi_n9_clk = clk;
	assign phi_n9_rst = rst;
	assign fork_24_in1_data = phi_n9_out1_data;
	assign fork_24_in1_valid = phi_n9_out1_valid;
	assign phi_n9_out1_ready = fork_24_in1_ready;

	assign fork_1_clk = clk;
	assign fork_1_rst = rst;
	assign add_13_in2_data = fork_1_out1_data;
	assign add_13_in2_valid = fork_1_out1_valid;
	assign fork_1_out1_ready = add_13_in2_ready;
	assign shl_17_in1_data = fork_1_out2_data;
	assign shl_17_in1_valid = fork_1_out2_valid;
	assign fork_1_out2_ready = shl_17_in1_ready;
	assign add_24_in1_data = fork_1_out3_data;
	assign add_24_in1_valid = fork_1_out3_valid;
	assign fork_1_out3_ready = add_24_in1_ready;

	assign fork_3_clk = clk;
	assign fork_3_rst = rst;
	assign icmp_25_in1_data = fork_3_out1_data;
	assign icmp_25_in1_valid = fork_3_out1_valid;
	assign fork_3_out1_ready = icmp_25_in1_ready;
	assign branch_8_in1_data = fork_3_out2_data;
	assign branch_8_in1_valid = fork_3_out2_valid;
	assign fork_3_out2_ready = branch_8_in1_ready;

	assign fork_23_clk = clk;
	assign fork_23_rst = rst;
	assign shl_12_in1_data = fork_23_out1_data;
	assign shl_12_in1_valid = fork_23_out1_valid;
	assign fork_23_out1_ready = shl_12_in1_ready;
	assign branch_9_in1_data = fork_23_out2_data;
	assign branch_9_in1_valid = fork_23_out2_valid;
	assign fork_23_out2_ready = branch_9_in1_ready;

	assign fork_24_clk = clk;
	assign fork_24_rst = rst;
	assign add_18_in2_data = fork_24_out1_data;
	assign add_18_in2_valid = fork_24_out1_valid;
	assign fork_24_out1_ready = add_18_in2_ready;
	assign branch_10_in1_data = fork_24_out2_data;
	assign branch_10_in1_valid = fork_24_out2_valid;
	assign fork_24_out2_ready = branch_10_in1_ready;

	assign branch_7_clk = clk;
	assign branch_7_rst = rst;
	assign Buffer_100_in1_data = branch_7_out1_data;
	assign Buffer_100_in1_valid = branch_7_out1_valid;
	assign branch_7_out1_ready = Buffer_100_in1_ready;
	assign phi_n7_in1_data = branch_7_out2_data;
	assign phi_n7_in1_valid = branch_7_out2_valid;
	assign branch_7_out2_ready = phi_n7_in1_ready;

	assign branch_8_clk = clk;
	assign branch_8_rst = rst;
	assign Buffer_101_in1_data = branch_8_out1_data;
	assign Buffer_101_in1_valid = branch_8_out1_valid;
	assign branch_8_out1_ready = Buffer_101_in1_ready;
	assign sink_7_in1_data = branch_8_out2_data;
	assign sink_7_in1_valid = branch_8_out2_valid;
	assign branch_8_out2_ready = sink_7_in1_ready;

	assign branch_9_clk = clk;
	assign branch_9_rst = rst;
	assign Buffer_102_in1_data = branch_9_out1_data;
	assign Buffer_102_in1_valid = branch_9_out1_valid;
	assign branch_9_out1_ready = Buffer_102_in1_ready;
	assign phi_n5_in1_data = branch_9_out2_data;
	assign phi_n5_in1_valid = branch_9_out2_valid;
	assign branch_9_out2_ready = phi_n5_in1_ready;

	assign branch_10_clk = clk;
	assign branch_10_rst = rst;
	assign Buffer_103_in1_data = branch_10_out1_data;
	assign Buffer_103_in1_valid = branch_10_out1_valid;
	assign branch_10_out1_ready = Buffer_103_in1_ready;
	assign phi_n6_in1_data = branch_10_out2_data;
	assign phi_n6_in1_valid = branch_10_out2_valid;
	assign branch_10_out2_ready = phi_n6_in1_ready;

	assign fork_36_clk = clk;
	assign fork_36_rst = rst;
	assign branch_10_in2_data = fork_36_out1_data;
	assign branch_10_in2_valid = fork_36_out1_valid;
	assign fork_36_out1_ready = branch_10_in2_ready;
	assign branch_9_in2_data = fork_36_out2_data;
	assign branch_9_in2_valid = fork_36_out2_valid;
	assign fork_36_out2_ready = branch_9_in2_ready;
	assign branch_8_in2_data = fork_36_out3_data;
	assign branch_8_in2_valid = fork_36_out3_valid;
	assign fork_36_out3_ready = branch_8_in2_ready;
	assign branch_7_in2_data = fork_36_out4_data;
	assign branch_7_in2_valid = fork_36_out4_valid;
	assign fork_36_out4_ready = branch_7_in2_ready;
	assign branchC_45_in2_data = fork_36_out5_data;
	assign branchC_45_in2_valid = fork_36_out5_valid;
	assign fork_36_out5_ready = branchC_45_in2_ready;

	assign phiC_23_clk = clk;
	assign phiC_23_rst = rst;
	assign branchC_45_in1_data = phiC_23_out1_data;
	assign branchC_45_in1_valid = phiC_23_out1_valid;
	assign phiC_23_out1_ready = branchC_45_in1_ready;
	assign fork_79_in1_data = phiC_23_out2_data;
	assign fork_79_in1_valid = phiC_23_out2_valid;
	assign phiC_23_out2_ready = fork_79_in1_ready;

	assign branchC_45_clk = clk;
	assign branchC_45_rst = rst;
	assign Buffer_104_in1_data = branchC_45_out1_data;
	assign Buffer_104_in1_valid = branchC_45_out1_valid;
	assign branchC_45_out1_ready = Buffer_104_in1_ready;
	assign phiC_24_in1_data = branchC_45_out2_data;
	assign phiC_24_in1_valid = branchC_45_out2_valid;
	assign branchC_45_out2_ready = phiC_24_in1_ready;

	assign source_1_clk = clk;
	assign source_1_rst = rst;
	assign cst_4_in1_data = source_1_out1_data;
	assign cst_4_in1_valid = source_1_out1_valid;
	assign source_1_out1_ready = cst_4_in1_ready;

	assign source_2_clk = clk;
	assign source_2_rst = rst;
	assign cst_5_in1_data = source_2_out1_data;
	assign cst_5_in1_valid = source_2_out1_valid;
	assign source_2_out1_ready = cst_5_in1_ready;

	assign source_3_clk = clk;
	assign source_3_rst = rst;
	assign cst_6_in1_data = source_3_out1_data;
	assign cst_6_in1_valid = source_3_out1_valid;
	assign source_3_out1_ready = cst_6_in1_ready;

	assign source_4_clk = clk;
	assign source_4_rst = rst;
	assign cst_7_in1_data = source_4_out1_data;
	assign cst_7_in1_valid = source_4_out1_valid;
	assign source_4_out1_ready = cst_7_in1_ready;

	assign fork_79_clk = clk;
	assign fork_79_rst = rst;
	assign phi_10_in1_data = fork_79_out1_data;
	assign phi_10_in1_valid = fork_79_out1_valid;
	assign fork_79_out1_ready = phi_10_in1_ready;
	assign phi_11_in1_data = fork_79_out2_data;
	assign phi_11_in1_valid = fork_79_out2_valid;
	assign fork_79_out2_ready = phi_11_in1_ready;

	assign phi_84_clk = clk;
	assign phi_84_rst = rst;
	assign and_305_in1_data = phi_84_out1_data;
	assign and_305_in1_valid = phi_84_out1_valid;
	assign phi_84_out1_ready = and_305_in1_ready;

	assign phi_85_clk = clk;
	assign phi_85_rst = rst;
	assign fork_13_in1_data = phi_85_out1_data;
	assign fork_13_in1_valid = phi_85_out1_valid;
	assign phi_85_out1_ready = fork_13_in1_ready;

	assign cst_30_clk = clk;
	assign cst_30_rst = rst;
	assign shl_86_in2_data = cst_30_out1_data;
	assign shl_86_in2_valid = cst_30_out1_valid;
	assign cst_30_out1_ready = shl_86_in2_ready;

	assign shl_86_clk = clk;
	assign shl_86_rst = rst;
	assign add_87_in1_data = shl_86_out1_data;
	assign add_87_in1_valid = shl_86_out1_valid;
	assign shl_86_out1_ready = add_87_in1_ready;

	assign add_87_clk = clk;
	assign add_87_rst = rst;
	assign load_90_in2_data = add_87_out1_data;
	assign load_90_in2_valid = add_87_out1_valid;
	assign add_87_out1_ready = load_90_in2_ready;

	assign load_90_clk = clk;
	assign load_90_rst = rst;
	assign and_304_in1_data = load_90_out1_data;
	assign and_304_in1_valid = load_90_out1_valid;
	assign load_90_out1_ready = and_304_in1_ready;
	assign MC_E_in5_data = load_90_out2_data;
	assign MC_E_in5_valid = load_90_out2_valid;
	assign load_90_out2_ready = MC_E_in5_ready;

	assign cst_31_clk = clk;
	assign cst_31_rst = rst;
	assign shl_91_in2_data = cst_31_out1_data;
	assign shl_91_in2_valid = cst_31_out1_valid;
	assign cst_31_out1_ready = shl_91_in2_ready;

	assign shl_91_clk = clk;
	assign shl_91_rst = rst;
	assign add_92_in1_data = shl_91_out1_data;
	assign add_92_in1_valid = shl_91_out1_valid;
	assign shl_91_out1_ready = add_92_in1_ready;

	assign add_92_clk = clk;
	assign add_92_rst = rst;
	assign load_95_in2_data = add_92_out1_data;
	assign load_95_in2_valid = add_92_out1_valid;
	assign add_92_out1_ready = load_95_in2_ready;

	assign load_95_clk = clk;
	assign load_95_rst = rst;
	assign and_304_in2_data = load_95_out1_data;
	assign and_304_in2_valid = load_95_out1_valid;
	assign load_95_out1_ready = and_304_in2_ready;
	assign MC_F_in5_data = load_95_out2_data;
	assign MC_F_in5_valid = load_95_out2_valid;
	assign load_95_out2_ready = MC_F_in5_ready;

	assign cst_32_clk = clk;
	assign cst_32_rst = rst;
	assign add_98_in2_data = cst_32_out1_data;
	assign add_98_in2_valid = cst_32_out1_valid;
	assign cst_32_out1_ready = add_98_in2_ready;

	assign add_98_clk = clk;
	assign add_98_rst = rst;
	assign fork_15_in1_data = add_98_out1_data;
	assign fork_15_in1_valid = add_98_out1_valid;
	assign add_98_out1_ready = fork_15_in1_ready;

	assign cst_33_clk = clk;
	assign cst_33_rst = rst;
	assign icmp_99_in2_data = cst_33_out1_data;
	assign icmp_99_in2_valid = cst_33_out1_valid;
	assign cst_33_out1_ready = icmp_99_in2_ready;

	assign icmp_99_clk = clk;
	assign icmp_99_rst = rst;
	assign fork_48_in1_data = icmp_99_out1_data;
	assign fork_48_in1_valid = icmp_99_out1_valid;
	assign icmp_99_out1_ready = fork_48_in1_ready;

	assign phi_n19_clk = clk;
	assign phi_n19_rst = rst;
	assign fork_31_in1_data = phi_n19_out1_data;
	assign fork_31_in1_valid = phi_n19_out1_valid;
	assign phi_n19_out1_ready = fork_31_in1_ready;

	assign phi_n20_clk = clk;
	assign phi_n20_rst = rst;
	assign fork_32_in1_data = phi_n20_out1_data;
	assign fork_32_in1_valid = phi_n20_out1_valid;
	assign phi_n20_out1_ready = fork_32_in1_ready;

	assign fork_13_clk = clk;
	assign fork_13_rst = rst;
	assign add_87_in2_data = fork_13_out1_data;
	assign add_87_in2_valid = fork_13_out1_valid;
	assign fork_13_out1_ready = add_87_in2_ready;
	assign shl_91_in1_data = fork_13_out2_data;
	assign shl_91_in1_valid = fork_13_out2_valid;
	assign fork_13_out2_ready = shl_91_in1_ready;
	assign add_98_in1_data = fork_13_out3_data;
	assign add_98_in1_valid = fork_13_out3_valid;
	assign fork_13_out3_ready = add_98_in1_ready;

	assign fork_15_clk = clk;
	assign fork_15_rst = rst;
	assign icmp_99_in1_data = fork_15_out1_data;
	assign icmp_99_in1_valid = fork_15_out1_valid;
	assign fork_15_out1_ready = icmp_99_in1_ready;
	assign branch_36_in1_data = fork_15_out2_data;
	assign branch_36_in1_valid = fork_15_out2_valid;
	assign fork_15_out2_ready = branch_36_in1_ready;

	assign fork_31_clk = clk;
	assign fork_31_rst = rst;
	assign shl_86_in1_data = fork_31_out1_data;
	assign shl_86_in1_valid = fork_31_out1_valid;
	assign fork_31_out1_ready = shl_86_in1_ready;
	assign branch_37_in1_data = fork_31_out2_data;
	assign branch_37_in1_valid = fork_31_out2_valid;
	assign fork_31_out2_ready = branch_37_in1_ready;

	assign fork_32_clk = clk;
	assign fork_32_rst = rst;
	assign add_92_in2_data = fork_32_out1_data;
	assign add_92_in2_valid = fork_32_out1_valid;
	assign fork_32_out1_ready = add_92_in2_ready;
	assign branch_38_in1_data = fork_32_out2_data;
	assign branch_38_in1_valid = fork_32_out2_valid;
	assign fork_32_out2_ready = branch_38_in1_ready;

	assign branch_35_clk = clk;
	assign branch_35_rst = rst;
	assign Buffer_120_in1_data = branch_35_out1_data;
	assign Buffer_120_in1_valid = branch_35_out1_valid;
	assign branch_35_out1_ready = Buffer_120_in1_ready;
	assign phi_n18_in1_data = branch_35_out2_data;
	assign phi_n18_in1_valid = branch_35_out2_valid;
	assign branch_35_out2_ready = phi_n18_in1_ready;

	assign branch_36_clk = clk;
	assign branch_36_rst = rst;
	assign Buffer_121_in1_data = branch_36_out1_data;
	assign Buffer_121_in1_valid = branch_36_out1_valid;
	assign branch_36_out1_ready = Buffer_121_in1_ready;
	assign sink_27_in1_data = branch_36_out2_data;
	assign sink_27_in1_valid = branch_36_out2_valid;
	assign branch_36_out2_ready = sink_27_in1_ready;

	assign branch_37_clk = clk;
	assign branch_37_rst = rst;
	assign Buffer_122_in1_data = branch_37_out1_data;
	assign Buffer_122_in1_valid = branch_37_out1_valid;
	assign branch_37_out1_ready = Buffer_122_in1_ready;
	assign phi_n16_in1_data = branch_37_out2_data;
	assign phi_n16_in1_valid = branch_37_out2_valid;
	assign branch_37_out2_ready = phi_n16_in1_ready;

	assign branch_38_clk = clk;
	assign branch_38_rst = rst;
	assign Buffer_123_in1_data = branch_38_out1_data;
	assign Buffer_123_in1_valid = branch_38_out1_valid;
	assign branch_38_out1_ready = Buffer_123_in1_ready;
	assign phi_n17_in1_data = branch_38_out2_data;
	assign phi_n17_in1_valid = branch_38_out2_valid;
	assign branch_38_out2_ready = phi_n17_in1_ready;

	assign fork_48_clk = clk;
	assign fork_48_rst = rst;
	assign branch_38_in2_data = fork_48_out1_data;
	assign branch_38_in2_valid = fork_48_out1_valid;
	assign fork_48_out1_ready = branch_38_in2_ready;
	assign branch_37_in2_data = fork_48_out2_data;
	assign branch_37_in2_valid = fork_48_out2_valid;
	assign fork_48_out2_ready = branch_37_in2_ready;
	assign branch_36_in2_data = fork_48_out3_data;
	assign branch_36_in2_valid = fork_48_out3_valid;
	assign fork_48_out3_ready = branch_36_in2_ready;
	assign branch_35_in2_data = fork_48_out4_data;
	assign branch_35_in2_valid = fork_48_out4_valid;
	assign fork_48_out4_ready = branch_35_in2_ready;
	assign branchC_57_in2_data = fork_48_out5_data;
	assign branchC_57_in2_valid = fork_48_out5_valid;
	assign fork_48_out5_ready = branchC_57_in2_ready;

	assign phiC_35_clk = clk;
	assign phiC_35_rst = rst;
	assign branchC_57_in1_data = phiC_35_out1_data;
	assign branchC_57_in1_valid = phiC_35_out1_valid;
	assign phiC_35_out1_ready = branchC_57_in1_ready;
	assign fork_85_in1_data = phiC_35_out2_data;
	assign fork_85_in1_valid = phiC_35_out2_valid;
	assign phiC_35_out2_ready = fork_85_in1_ready;

	assign branchC_57_clk = clk;
	assign branchC_57_rst = rst;
	assign Buffer_124_in1_data = branchC_57_out1_data;
	assign Buffer_124_in1_valid = branchC_57_out1_valid;
	assign branchC_57_out1_ready = Buffer_124_in1_ready;
	assign phiC_36_in1_data = branchC_57_out2_data;
	assign phiC_36_in1_valid = branchC_57_out2_valid;
	assign branchC_57_out2_ready = phiC_36_in1_ready;

	assign source_21_clk = clk;
	assign source_21_rst = rst;
	assign cst_30_in1_data = source_21_out1_data;
	assign cst_30_in1_valid = source_21_out1_valid;
	assign source_21_out1_ready = cst_30_in1_ready;

	assign source_22_clk = clk;
	assign source_22_rst = rst;
	assign cst_31_in1_data = source_22_out1_data;
	assign cst_31_in1_valid = source_22_out1_valid;
	assign source_22_out1_ready = cst_31_in1_ready;

	assign source_23_clk = clk;
	assign source_23_rst = rst;
	assign cst_32_in1_data = source_23_out1_data;
	assign cst_32_in1_valid = source_23_out1_valid;
	assign source_23_out1_ready = cst_32_in1_ready;

	assign source_24_clk = clk;
	assign source_24_rst = rst;
	assign cst_33_in1_data = source_24_out1_data;
	assign cst_33_in1_valid = source_24_out1_valid;
	assign source_24_out1_ready = cst_33_in1_ready;

	assign fork_85_clk = clk;
	assign fork_85_rst = rst;
	assign phi_84_in1_data = fork_85_out1_data;
	assign phi_84_in1_valid = fork_85_out1_valid;
	assign fork_85_out1_ready = phi_84_in1_ready;
	assign phi_85_in1_data = fork_85_out2_data;
	assign phi_85_in1_valid = fork_85_out2_valid;
	assign fork_85_out2_ready = phi_85_in1_ready;

	assign phi_1_clk = clk;
	assign phi_1_rst = rst;
	assign branch_2_in1_data = phi_1_out1_data;
	assign branch_2_in1_valid = phi_1_out1_valid;
	assign phi_1_out1_ready = branch_2_in1_ready;

	assign brCst_block2_clk = clk;
	assign brCst_block2_rst = rst;
	assign fork_34_in1_data = brCst_block2_out1_data;
	assign fork_34_in1_valid = brCst_block2_out1_valid;
	assign brCst_block2_out1_ready = fork_34_in1_ready;

	assign cst_1_clk = clk;
	assign cst_1_rst = rst;
	assign branch_1_in1_data = cst_1_out1_data;
	assign branch_1_in1_valid = cst_1_out1_valid;
	assign cst_1_out1_ready = branch_1_in1_ready;

	assign branch_1_clk = clk;
	assign branch_1_rst = rst;
	assign phi_3_in2_data = branch_1_out1_data;
	assign phi_3_in2_valid = branch_1_out1_valid;
	assign branch_1_out1_ready = phi_3_in2_ready;
	assign sink_1_in1_data = branch_1_out2_data;
	assign sink_1_in1_valid = branch_1_out2_valid;
	assign branch_1_out2_ready = sink_1_in1_ready;

	assign branch_2_clk = clk;
	assign branch_2_rst = rst;
	assign phi_n4_in1_data = branch_2_out1_data;
	assign phi_n4_in1_valid = branch_2_out1_valid;
	assign branch_2_out1_ready = phi_n4_in1_ready;
	assign sink_2_in1_data = branch_2_out2_data;
	assign sink_2_in1_valid = branch_2_out2_valid;
	assign branch_2_out2_ready = sink_2_in1_ready;

	assign fork_34_clk = clk;
	assign fork_34_rst = rst;
	assign branch_2_in2_data = fork_34_out1_data;
	assign branch_2_in2_valid = fork_34_out1_valid;
	assign fork_34_out1_ready = branch_2_in2_ready;
	assign branch_1_in2_data = fork_34_out2_data;
	assign branch_1_in2_valid = fork_34_out2_valid;
	assign fork_34_out2_ready = branch_1_in2_ready;
	assign branchC_43_in2_data = fork_34_out3_data;
	assign branchC_43_in2_valid = fork_34_out3_valid;
	assign fork_34_out3_ready = branchC_43_in2_ready;

	assign phiC_21_clk = clk;
	assign phiC_21_rst = rst;
	assign forkC_54_in1_data = phiC_21_out1_data;
	assign forkC_54_in1_valid = phiC_21_out1_valid;
	assign phiC_21_out1_ready = forkC_54_in1_ready;
	assign phi_1_in1_data = phiC_21_out2_data;
	assign phi_1_in1_valid = phiC_21_out2_valid;
	assign phiC_21_out2_ready = phi_1_in1_ready;

	assign forkC_54_clk = clk;
	assign forkC_54_rst = rst;
	assign cst_1_in1_data = forkC_54_out1_data;
	assign cst_1_in1_valid = forkC_54_out1_valid;
	assign forkC_54_out1_ready = cst_1_in1_ready;
	assign branchC_43_in1_data = forkC_54_out2_data;
	assign branchC_43_in1_valid = forkC_54_out2_valid;
	assign forkC_54_out2_ready = branchC_43_in1_ready;
	assign brCst_block2_in1_data = forkC_54_out3_data;
	assign brCst_block2_in1_valid = forkC_54_out3_valid;
	assign forkC_54_out3_ready = brCst_block2_in1_ready;

	assign branchC_43_clk = clk;
	assign branchC_43_rst = rst;
	assign phiC_22_in1_data = branchC_43_out1_data;
	assign phiC_22_in1_valid = branchC_43_out1_valid;
	assign branchC_43_out1_ready = phiC_22_in1_ready;
	assign sink_31_in1_data = branchC_43_out2_data;
	assign sink_31_in1_valid = branchC_43_out2_valid;
	assign branchC_43_out2_ready = sink_31_in1_ready;

	assign MC_E_clk = clk;
	assign MC_E_rst = rst;
	assign E_ce0 = E_we0;
	assign load_8_in1_data = MC_E_out1_data;
	assign load_8_in1_valid = MC_E_out1_valid;
	assign MC_E_out1_ready = load_8_in1_ready;
	assign load_90_in1_data = MC_E_out2_data;
	assign load_90_in1_valid = MC_E_out2_valid;
	assign MC_E_out2_ready = load_90_in1_ready;
	assign end_0_in1_data = MC_E_out3_data;
	assign end_0_in1_valid = MC_E_out3_valid;
	assign MC_E_out3_ready = end_0_in1_ready;

	assign MC_A_clk = clk;
	assign MC_A_rst = rst;
	assign A_ce0 = A_we0;
	assign MC_A_in2_valid = 0;
	assign MC_A_in2_data = 0;
	assign load_16_in1_data = MC_A_out1_data;
	assign load_16_in1_valid = MC_A_out1_valid;
	assign MC_A_out1_ready = load_16_in1_ready;
	assign end_0_in2_data = MC_A_out2_data;
	assign end_0_in2_valid = MC_A_out2_valid;
	assign MC_A_out2_ready = end_0_in2_ready;

	assign MC_B_clk = clk;
	assign MC_B_rst = rst;
	assign B_ce0 = B_we0;
	assign MC_B_in2_valid = 0;
	assign MC_B_in2_data = 0;
	assign load_21_in1_data = MC_B_out1_data;
	assign load_21_in1_valid = MC_B_out1_valid;
	assign MC_B_out1_ready = load_21_in1_ready;
	assign end_0_in3_data = MC_B_out2_data;
	assign end_0_in3_valid = MC_B_out2_valid;
	assign MC_B_out2_ready = end_0_in3_ready;

	assign MC_F_clk = clk;
	assign MC_F_rst = rst;
	assign F_ce0 = F_we0;
	assign load_45_in1_data = MC_F_out1_data;
	assign load_45_in1_valid = MC_F_out1_valid;
	assign MC_F_out1_ready = load_45_in1_ready;
	assign load_95_in1_data = MC_F_out2_data;
	assign load_95_in1_valid = MC_F_out2_valid;
	assign MC_F_out2_ready = load_95_in1_ready;
	assign end_0_in4_data = MC_F_out3_data;
	assign end_0_in4_valid = MC_F_out3_valid;
	assign MC_F_out3_ready = end_0_in4_ready;

	assign MC_C_clk = clk;
	assign MC_C_rst = rst;
	assign C_ce0 = C_we0;
	assign MC_C_in2_valid = 0;
	assign MC_C_in2_data = 0;
	assign load_53_in1_data = MC_C_out1_data;
	assign load_53_in1_valid = MC_C_out1_valid;
	assign MC_C_out1_ready = load_53_in1_ready;
	assign end_0_in5_data = MC_C_out2_data;
	assign end_0_in5_valid = MC_C_out2_valid;
	assign MC_C_out2_ready = end_0_in5_ready;

	assign MC_D_clk = clk;
	assign MC_D_rst = rst;
	assign D_ce0 = D_we0;
	assign MC_D_in2_valid = 0;
	assign MC_D_in2_data = 0;
	assign load_58_in1_data = MC_D_out1_data;
	assign load_58_in1_valid = MC_D_out1_valid;
	assign MC_D_out1_ready = load_58_in1_ready;
	assign end_0_in6_data = MC_D_out2_data;
	assign end_0_in6_valid = MC_D_out2_valid;
	assign MC_D_out2_ready = end_0_in6_ready;

	assign MC_G_clk = clk;
	assign MC_G_rst = rst;
	assign G_ce0 = G_we0;
	assign load_82_in1_data = MC_G_out1_data;
	assign load_82_in1_valid = MC_G_out1_valid;
	assign MC_G_out1_ready = load_82_in1_ready;
	assign end_0_in7_data = MC_G_out2_data;
	assign end_0_in7_valid = MC_G_out2_valid;
	assign MC_G_out2_ready = end_0_in7_ready;

	assign sink_0_clk = clk;
	assign sink_0_rst = rst;

	assign sink_1_clk = clk;
	assign sink_1_rst = rst;

	assign sink_2_clk = clk;
	assign sink_2_rst = rst;

	assign sink_3_clk = clk;
	assign sink_3_rst = rst;

	assign sink_4_clk = clk;
	assign sink_4_rst = rst;

	assign sink_5_clk = clk;
	assign sink_5_rst = rst;

	assign sink_6_clk = clk;
	assign sink_6_rst = rst;

	assign sink_7_clk = clk;
	assign sink_7_rst = rst;

	assign sink_8_clk = clk;
	assign sink_8_rst = rst;

	assign sink_9_clk = clk;
	assign sink_9_rst = rst;

	assign sink_10_clk = clk;
	assign sink_10_rst = rst;

	assign sink_11_clk = clk;
	assign sink_11_rst = rst;

	assign sink_12_clk = clk;
	assign sink_12_rst = rst;

	assign sink_13_clk = clk;
	assign sink_13_rst = rst;

	assign sink_14_clk = clk;
	assign sink_14_rst = rst;

	assign sink_15_clk = clk;
	assign sink_15_rst = rst;

	assign sink_16_clk = clk;
	assign sink_16_rst = rst;

	assign sink_17_clk = clk;
	assign sink_17_rst = rst;

	assign sink_18_clk = clk;
	assign sink_18_rst = rst;

	assign sink_19_clk = clk;
	assign sink_19_rst = rst;

	assign sink_20_clk = clk;
	assign sink_20_rst = rst;

	assign sink_21_clk = clk;
	assign sink_21_rst = rst;

	assign sink_22_clk = clk;
	assign sink_22_rst = rst;

	assign sink_23_clk = clk;
	assign sink_23_rst = rst;

	assign sink_24_clk = clk;
	assign sink_24_rst = rst;

	assign sink_25_clk = clk;
	assign sink_25_rst = rst;

	assign sink_26_clk = clk;
	assign sink_26_rst = rst;

	assign sink_27_clk = clk;
	assign sink_27_rst = rst;

	assign sink_28_clk = clk;
	assign sink_28_rst = rst;

	assign sink_29_clk = clk;
	assign sink_29_rst = rst;

	assign sink_30_clk = clk;
	assign sink_30_rst = rst;

	assign sink_31_clk = clk;
	assign sink_31_rst = rst;

	assign sink_32_clk = clk;
	assign sink_32_rst = rst;

	assign sink_33_clk = clk;
	assign sink_33_rst = rst;

	assign sink_34_clk = clk;
	assign sink_34_rst = rst;

	assign sink_35_clk = clk;
	assign sink_35_rst = rst;

	assign sink_36_clk = clk;
	assign sink_36_rst = rst;

	assign sink_37_clk = clk;
	assign sink_37_rst = rst;

	assign sink_38_clk = clk;
	assign sink_38_rst = rst;

	assign Buffer_100_clk = clk;
	assign Buffer_100_rst = rst;
	assign phi_10_in3_data = Buffer_100_out1_data;
	assign phi_10_in3_valid = Buffer_100_out1_valid;
	assign Buffer_100_out1_ready = phi_10_in3_ready;

	assign Buffer_101_clk = clk;
	assign Buffer_101_rst = rst;
	assign phi_11_in3_data = Buffer_101_out1_data;
	assign phi_11_in3_valid = Buffer_101_out1_valid;
	assign Buffer_101_out1_ready = phi_11_in3_ready;

	assign Buffer_102_clk = clk;
	assign Buffer_102_rst = rst;
	assign phi_n8_in2_data = Buffer_102_out1_data;
	assign phi_n8_in2_valid = Buffer_102_out1_valid;
	assign Buffer_102_out1_ready = phi_n8_in2_ready;

	assign Buffer_103_clk = clk;
	assign Buffer_103_rst = rst;
	assign phi_n9_in2_data = Buffer_103_out1_data;
	assign phi_n9_in2_valid = Buffer_103_out1_valid;
	assign Buffer_103_out1_ready = phi_n9_in2_ready;

	assign Buffer_104_clk = clk;
	assign Buffer_104_rst = rst;
	assign phiC_23_in2_data = Buffer_104_out1_data;
	assign phiC_23_in2_valid = Buffer_104_out1_valid;
	assign Buffer_104_out1_ready = phiC_23_in2_ready;

	assign Buffer_105_clk = clk;
	assign Buffer_105_rst = rst;
	assign phi_3_in3_data = Buffer_105_out1_data;
	assign phi_3_in3_valid = Buffer_105_out1_valid;
	assign Buffer_105_out1_ready = phi_3_in3_ready;

	assign Buffer_106_clk = clk;
	assign Buffer_106_rst = rst;
	assign phi_n4_in2_data = Buffer_106_out1_data;
	assign phi_n4_in2_valid = Buffer_106_out1_valid;
	assign Buffer_106_out1_ready = phi_n4_in2_ready;

	assign Buffer_107_clk = clk;
	assign Buffer_107_rst = rst;
	assign phiC_22_in2_data = Buffer_107_out1_data;
	assign phiC_22_in2_valid = Buffer_107_out1_valid;
	assign Buffer_107_out1_ready = phiC_22_in2_ready;

	assign Buffer_108_clk = clk;
	assign Buffer_108_rst = rst;
	assign phi_1_in3_data = Buffer_108_out1_data;
	assign phi_1_in3_valid = Buffer_108_out1_valid;
	assign Buffer_108_out1_ready = phi_1_in3_ready;

	assign Buffer_109_clk = clk;
	assign Buffer_109_rst = rst;
	assign phiC_21_in2_data = Buffer_109_out1_data;
	assign phiC_21_in2_valid = Buffer_109_out1_valid;
	assign Buffer_109_out1_ready = phiC_21_in2_ready;

	assign Buffer_110_clk = clk;
	assign Buffer_110_rst = rst;
	assign phi_47_in3_data = Buffer_110_out1_data;
	assign phi_47_in3_valid = Buffer_110_out1_valid;
	assign Buffer_110_out1_ready = phi_47_in3_ready;

	assign Buffer_111_clk = clk;
	assign Buffer_111_rst = rst;
	assign phi_48_in3_data = Buffer_111_out1_data;
	assign phi_48_in3_valid = Buffer_111_out1_valid;
	assign Buffer_111_out1_ready = phi_48_in3_ready;

	assign Buffer_112_clk = clk;
	assign Buffer_112_rst = rst;
	assign phi_n10_in2_data = Buffer_112_out1_data;
	assign phi_n10_in2_valid = Buffer_112_out1_valid;
	assign Buffer_112_out1_ready = phi_n10_in2_ready;

	assign Buffer_113_clk = clk;
	assign Buffer_113_rst = rst;
	assign phi_n11_in2_data = Buffer_113_out1_data;
	assign phi_n11_in2_valid = Buffer_113_out1_valid;
	assign Buffer_113_out1_ready = phi_n11_in2_ready;

	assign Buffer_114_clk = clk;
	assign Buffer_114_rst = rst;
	assign phiC_29_in2_data = Buffer_114_out1_data;
	assign phiC_29_in2_valid = Buffer_114_out1_valid;
	assign Buffer_114_out1_ready = phiC_29_in2_ready;

	assign Buffer_115_clk = clk;
	assign Buffer_115_rst = rst;
	assign phi_40_in3_data = Buffer_115_out1_data;
	assign phi_40_in3_valid = Buffer_115_out1_valid;
	assign Buffer_115_out1_ready = phi_40_in3_ready;

	assign Buffer_116_clk = clk;
	assign Buffer_116_rst = rst;
	assign phi_n13_in2_data = Buffer_116_out1_data;
	assign phi_n13_in2_valid = Buffer_116_out1_valid;
	assign Buffer_116_out1_ready = phi_n13_in2_ready;

	assign Buffer_117_clk = clk;
	assign Buffer_117_rst = rst;
	assign phiC_28_in2_data = Buffer_117_out1_data;
	assign phiC_28_in2_valid = Buffer_117_out1_valid;
	assign Buffer_117_out1_ready = phiC_28_in2_ready;

	assign Buffer_118_clk = clk;
	assign Buffer_118_rst = rst;
	assign phi_38_in3_data = Buffer_118_out1_data;
	assign phi_38_in3_valid = Buffer_118_out1_valid;
	assign Buffer_118_out1_ready = phi_38_in3_ready;

	assign Buffer_119_clk = clk;
	assign Buffer_119_rst = rst;
	assign phiC_27_in2_data = Buffer_119_out1_data;
	assign phiC_27_in2_valid = Buffer_119_out1_valid;
	assign Buffer_119_out1_ready = phiC_27_in2_ready;

	assign Buffer_120_clk = clk;
	assign Buffer_120_rst = rst;
	assign phi_84_in3_data = Buffer_120_out1_data;
	assign phi_84_in3_valid = Buffer_120_out1_valid;
	assign Buffer_120_out1_ready = phi_84_in3_ready;

	assign Buffer_121_clk = clk;
	assign Buffer_121_rst = rst;
	assign phi_85_in3_data = Buffer_121_out1_data;
	assign phi_85_in3_valid = Buffer_121_out1_valid;
	assign Buffer_121_out1_ready = phi_85_in3_ready;

	assign Buffer_122_clk = clk;
	assign Buffer_122_rst = rst;
	assign phi_n19_in2_data = Buffer_122_out1_data;
	assign phi_n19_in2_valid = Buffer_122_out1_valid;
	assign Buffer_122_out1_ready = phi_n19_in2_ready;

	assign Buffer_123_clk = clk;
	assign Buffer_123_rst = rst;
	assign phi_n20_in2_data = Buffer_123_out1_data;
	assign phi_n20_in2_valid = Buffer_123_out1_valid;
	assign Buffer_123_out1_ready = phi_n20_in2_ready;

	assign Buffer_124_clk = clk;
	assign Buffer_124_rst = rst;
	assign phiC_35_in2_data = Buffer_124_out1_data;
	assign phiC_35_in2_valid = Buffer_124_out1_valid;
	assign Buffer_124_out1_ready = phiC_35_in2_ready;

	assign Buffer_125_clk = clk;
	assign Buffer_125_rst = rst;
	assign phi_77_in3_data = Buffer_125_out1_data;
	assign phi_77_in3_valid = Buffer_125_out1_valid;
	assign Buffer_125_out1_ready = phi_77_in3_ready;

	assign Buffer_126_clk = clk;
	assign Buffer_126_rst = rst;
	assign phi_n15_in2_data = Buffer_126_out1_data;
	assign phi_n15_in2_valid = Buffer_126_out1_valid;
	assign Buffer_126_out1_ready = phi_n15_in2_ready;

	assign Buffer_127_clk = clk;
	assign Buffer_127_rst = rst;
	assign phiC_34_in2_data = Buffer_127_out1_data;
	assign phiC_34_in2_valid = Buffer_127_out1_valid;
	assign Buffer_127_out1_ready = phiC_34_in2_ready;

	assign Buffer_128_clk = clk;
	assign Buffer_128_rst = rst;
	assign phi_75_in3_data = Buffer_128_out1_data;
	assign phi_75_in3_valid = Buffer_128_out1_valid;
	assign Buffer_128_out1_ready = phi_75_in3_ready;

	assign Buffer_129_clk = clk;
	assign Buffer_129_rst = rst;
	assign phiC_33_in2_data = Buffer_129_out1_data;
	assign phiC_33_in2_valid = Buffer_129_out1_valid;
	assign Buffer_129_out1_ready = phiC_33_in2_ready;

	assign and_300_clk = clk;
	assign and_300_rst = rst;
	assign Buffer_300_in1_data = and_300_out1_data;
	assign Buffer_300_in1_valid = and_300_out1_valid;
	assign and_300_out1_ready = Buffer_300_in1_ready;

	assign Buffer_300_clk = clk;
	assign Buffer_300_rst = rst;
	assign and_301_in2_data = Buffer_300_out1_data;
	assign and_301_in2_valid = Buffer_300_out1_valid;
	assign Buffer_300_out1_ready = and_301_in2_ready;

	assign and_301_clk = clk;
	assign and_301_rst = rst;
	assign Buffer_301_in1_data = and_301_out1_data;
	assign Buffer_301_in1_valid = and_301_out1_valid;
	assign and_301_out1_ready = Buffer_301_in1_ready;

	assign Buffer_301_clk = clk;
	assign Buffer_301_rst = rst;
	assign branch_7_in1_data = Buffer_301_out1_data;
	assign branch_7_in1_valid = Buffer_301_out1_valid;
	assign Buffer_301_out1_ready = branch_7_in1_ready;

	assign and_302_clk = clk;
	assign and_302_rst = rst;
	assign Buffer_302_in1_data = and_302_out1_data;
	assign Buffer_302_in1_valid = and_302_out1_valid;
	assign and_302_out1_ready = Buffer_302_in1_ready;

	assign Buffer_302_clk = clk;
	assign Buffer_302_rst = rst;
	assign and_303_in2_data = Buffer_302_out1_data;
	assign and_303_in2_valid = Buffer_302_out1_valid;
	assign Buffer_302_out1_ready = and_303_in2_ready;

	assign and_303_clk = clk;
	assign and_303_rst = rst;
	assign Buffer_303_in1_data = and_303_out1_data;
	assign Buffer_303_in1_valid = and_303_out1_valid;
	assign and_303_out1_ready = Buffer_303_in1_ready;

	assign Buffer_303_clk = clk;
	assign Buffer_303_rst = rst;
	assign branch_21_in1_data = Buffer_303_out1_data;
	assign branch_21_in1_valid = Buffer_303_out1_valid;
	assign Buffer_303_out1_ready = branch_21_in1_ready;

	assign and_304_clk = clk;
	assign and_304_rst = rst;
	assign Buffer_304_in1_data = and_304_out1_data;
	assign Buffer_304_in1_valid = and_304_out1_valid;
	assign and_304_out1_ready = Buffer_304_in1_ready;

	assign Buffer_304_clk = clk;
	assign Buffer_304_rst = rst;
	assign and_305_in2_data = Buffer_304_out1_data;
	assign and_305_in2_valid = Buffer_304_out1_valid;
	assign Buffer_304_out1_ready = and_305_in2_ready;

	assign and_305_clk = clk;
	assign and_305_rst = rst;
	assign Buffer_305_in1_data = and_305_out1_data;
	assign Buffer_305_in1_valid = and_305_out1_valid;
	assign and_305_out1_ready = Buffer_305_in1_ready;

	assign Buffer_305_clk = clk;
	assign Buffer_305_rst = rst;
	assign branch_35_in1_data = Buffer_305_out1_data;
	assign branch_35_in1_valid = Buffer_305_out1_valid;
	assign Buffer_305_out1_ready = branch_35_in1_ready;

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4), .COND_SIZE(1)) mux_node_phi_3
		(.clk(phi_3_clk), .rst(phi_3_rst),
		.data_in_bus({{3'b0, phi_3_in1_data}, phi_3_in3_data, phi_3_in2_data}), .valid_in_bus({phi_3_in1_valid, phi_3_in3_valid, phi_3_in2_valid}), .ready_in_bus({phi_3_in1_ready, phi_3_in3_ready, phi_3_in2_ready}), 
		.data_out_bus({phi_3_out1_data}), .valid_out_bus({phi_3_out1_valid}), .ready_out_bus({phi_3_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_2
		(.clk(cst_2_clk), .rst(cst_2_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_2_in1_valid}), .ready_in_bus({cst_2_in1_ready}), 
		.data_out_bus({cst_2_out1_data}), .valid_out_bus({cst_2_out1_valid}), .ready_out_bus({cst_2_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_4
		(.clk(shl_4_clk), .rst(shl_4_rst),
		.data_in_bus({shl_4_in2_data, shl_4_in1_data}), .valid_in_bus({shl_4_in2_valid, shl_4_in1_valid}), .ready_in_bus({shl_4_in2_ready, shl_4_in1_ready}), 
		.data_out_bus({shl_4_out1_data}), .valid_out_bus({shl_4_out1_valid}), .ready_out_bus({shl_4_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_5
		(.clk(add_5_clk), .rst(add_5_rst),
		.data_in_bus({add_5_in2_data, add_5_in1_data}), .valid_in_bus({add_5_in2_valid, add_5_in1_valid}), .ready_in_bus({add_5_in2_ready, add_5_in1_ready}), 
		.data_out_bus({add_5_out1_data}), .valid_out_bus({add_5_out1_valid}), .ready_out_bus({add_5_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_load_op_load_8
		(.clk(load_8_clk), .rst(load_8_rst),
		.data_in_bus({load_8_in1_data}), .address_in_bus({load_8_in2_data}), .valid_in_bus({load_8_in2_valid, load_8_in1_valid}), .ready_in_bus({load_8_in2_ready, load_8_in1_ready}), 
		.data_out_bus({load_8_out1_data}), .address_out_bus({load_8_out2_data}), .valid_out_bus({load_8_out2_valid, load_8_out1_valid}), .ready_out_bus({load_8_out2_ready, load_8_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block3
		(.clk(brCst_block3_clk), .rst(brCst_block3_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block3_in1_valid}), .ready_in_bus({brCst_block3_in1_ready}), 
		.data_out_bus({brCst_block3_out1_data}), .valid_out_bus({brCst_block3_out1_valid}), .ready_out_bus({brCst_block3_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_3
		(.clk(cst_3_clk), .rst(cst_3_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_3_in1_valid}), .ready_in_bus({cst_3_in1_ready}), 
		.data_out_bus({cst_3_out1_data}), .valid_out_bus({cst_3_out1_valid}), .ready_out_bus({cst_3_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n4
		(.clk(phi_n4_clk), .rst(phi_n4_rst),
		.data_in_bus({phi_n4_in2_data, phi_n4_in1_data}), .valid_in_bus({phi_n4_in2_valid, phi_n4_in1_valid}), .ready_in_bus({phi_n4_in2_ready, phi_n4_in1_ready}), 
		.data_out_bus({phi_n4_out1_data}), .valid_out_bus({phi_n4_out1_valid}), .ready_out_bus({phi_n4_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_0
		(.clk(fork_0_clk), .rst(fork_0_rst),
		.data_in_bus({fork_0_in1_data}), .valid_in_bus({fork_0_in1_valid}), .ready_in_bus({fork_0_in1_ready}), 
		.data_out_bus({fork_0_out2_data, fork_0_out1_data}), .valid_out_bus({fork_0_out2_valid, fork_0_out1_valid}), .ready_out_bus({fork_0_out2_ready, fork_0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_20
		(.clk(fork_20_clk), .rst(fork_20_rst),
		.data_in_bus({fork_20_in1_data}), .valid_in_bus({fork_20_in1_valid}), .ready_in_bus({fork_20_in1_ready}), 
		.data_out_bus({fork_20_out2_data, fork_20_out1_data}), .valid_out_bus({fork_20_out2_valid, fork_20_out1_valid}), .ready_out_bus({fork_20_out2_ready, fork_20_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_3
		(.clk(branch_3_clk), .rst(branch_3_rst),
		.data_in_bus({{31'b0, branch_3_in2_data}, branch_3_in1_data}), .valid_in_bus({branch_3_in2_valid, branch_3_in1_valid}), .ready_in_bus({branch_3_in2_ready, branch_3_in1_ready}), 
		.data_out_bus({branch_3_out2_data, branch_3_out1_data}), .valid_out_bus({branch_3_out2_valid, branch_3_out1_valid}), .ready_out_bus({branch_3_out2_ready, branch_3_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_4
		(.clk(branch_4_clk), .rst(branch_4_rst),
		.data_in_bus({{branch_4_in2_data}, branch_4_in1_data}), .valid_in_bus({branch_4_in2_valid, branch_4_in1_valid}), .ready_in_bus({branch_4_in2_ready, branch_4_in1_ready}), 
		.data_out_bus({branch_4_out2_data, branch_4_out1_data}), .valid_out_bus({branch_4_out2_valid, branch_4_out1_valid}), .ready_out_bus({branch_4_out2_ready, branch_4_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_5
		(.clk(branch_5_clk), .rst(branch_5_rst),
		.data_in_bus({{3'b0, branch_5_in2_data}, branch_5_in1_data}), .valid_in_bus({branch_5_in2_valid, branch_5_in1_valid}), .ready_in_bus({branch_5_in2_ready, branch_5_in1_ready}), 
		.data_out_bus({branch_5_out2_data, branch_5_out1_data}), .valid_out_bus({branch_5_out2_valid, branch_5_out1_valid}), .ready_out_bus({branch_5_out2_ready, branch_5_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_6
		(.clk(branch_6_clk), .rst(branch_6_rst),
		.data_in_bus({{3'b0, branch_6_in2_data}, branch_6_in1_data}), .valid_in_bus({branch_6_in2_valid, branch_6_in1_valid}), .ready_in_bus({branch_6_in2_ready, branch_6_in1_ready}), 
		.data_out_bus({branch_6_out2_data, branch_6_out1_data}), .valid_out_bus({branch_6_out2_valid, branch_6_out1_valid}), .ready_out_bus({branch_6_out2_ready, branch_6_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_35
		(.clk(fork_35_clk), .rst(fork_35_rst),
		.data_in_bus({fork_35_in1_data}), .valid_in_bus({fork_35_in1_valid}), .ready_in_bus({fork_35_in1_ready}), 
		.data_out_bus({fork_35_out5_data, fork_35_out4_data, fork_35_out3_data, fork_35_out2_data, fork_35_out1_data}), .valid_out_bus({fork_35_out5_valid, fork_35_out4_valid, fork_35_out3_valid, fork_35_out2_valid, fork_35_out1_valid}), .ready_out_bus({fork_35_out5_ready, fork_35_out4_ready, fork_35_out3_ready, fork_35_out2_ready, fork_35_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_22
		(.clk(phiC_22_clk), .rst(phiC_22_rst),
		.data_in_bus({phiC_22_in2_data, phiC_22_in1_data}), .valid_in_bus({phiC_22_in2_valid, phiC_22_in1_valid}), .ready_in_bus({phiC_22_in2_ready, phiC_22_in1_ready}), 
		.data_out_bus({phiC_22_out2_data, phiC_22_out1_data}), .valid_out_bus({phiC_22_out2_valid, phiC_22_out1_valid}), .ready_out_bus({phiC_22_out2_ready, phiC_22_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_55
		(.clk(forkC_55_clk), .rst(forkC_55_rst),
		.data_in_bus({forkC_55_in1_data}), .valid_in_bus({forkC_55_in1_valid}), .ready_in_bus({forkC_55_in1_ready}), 
		.data_out_bus({forkC_55_out3_data, forkC_55_out2_data, forkC_55_out1_data}), .valid_out_bus({forkC_55_out3_valid, forkC_55_out2_valid, forkC_55_out1_valid}), .ready_out_bus({forkC_55_out3_ready, forkC_55_out2_ready, forkC_55_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_44
		(.clk(branchC_44_clk), .rst(branchC_44_rst),
		.data_in_bus({{branchC_44_in2_data}, branchC_44_in1_data}), .valid_in_bus({branchC_44_in2_valid, branchC_44_in1_valid}), .ready_in_bus({branchC_44_in2_ready, branchC_44_in1_ready}), 
		.data_out_bus({branchC_44_out2_data, branchC_44_out1_data}), .valid_out_bus({branchC_44_out2_valid, branchC_44_out1_valid}), .ready_out_bus({branchC_44_out2_ready, branchC_44_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_0
		(.clk(source_0_clk), .rst(source_0_rst),
		.data_out_bus({source_0_out1_data}), .valid_out_bus({source_0_out1_valid}), .ready_out_bus({source_0_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_8
		(.clk(cst_8_clk), .rst(cst_8_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_8_in1_valid}), .ready_in_bus({cst_8_in1_ready}), 
		.data_out_bus({cst_8_out1_data}), .valid_out_bus({cst_8_out1_valid}), .ready_out_bus({cst_8_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_27
		(.clk(shl_27_clk), .rst(shl_27_rst),
		.data_in_bus({shl_27_in2_data, shl_27_in1_data}), .valid_in_bus({shl_27_in2_valid, shl_27_in1_valid}), .ready_in_bus({shl_27_in2_ready, shl_27_in1_ready}), 
		.data_out_bus({shl_27_out1_data}), .valid_out_bus({shl_27_out1_valid}), .ready_out_bus({shl_27_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_28
		(.clk(add_28_clk), .rst(add_28_rst),
		.data_in_bus({add_28_in2_data, add_28_in1_data}), .valid_in_bus({add_28_in2_valid, add_28_in1_valid}), .ready_in_bus({add_28_in2_ready, add_28_in1_ready}), 
		.data_out_bus({add_28_out1_data}), .valid_out_bus({add_28_out1_valid}), .ready_out_bus({add_28_out1_ready}));

	mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_store_op_store_0
		(.clk(store_0_clk), .rst(store_0_rst),
		.data_in_bus({store_0_in1_data}), .address_in_bus({store_0_in2_data}), .valid_in_bus({store_0_in2_valid, store_0_in1_valid}), .ready_in_bus({store_0_in2_ready, store_0_in1_ready}), 
		.data_out_bus({store_0_out1_data}), .address_out_bus({store_0_out2_data}), .valid_out_bus({store_0_out2_valid, store_0_out1_valid}), .ready_out_bus({store_0_out2_ready, store_0_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_9
		(.clk(cst_9_clk), .rst(cst_9_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_9_in1_valid}), .ready_in_bus({cst_9_in1_ready}), 
		.data_out_bus({cst_9_out1_data}), .valid_out_bus({cst_9_out1_valid}), .ready_out_bus({cst_9_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) add_op_add_31
		(.clk(add_31_clk), .rst(add_31_rst),
		.data_in_bus({add_31_in2_data, add_31_in1_data}), .valid_in_bus({add_31_in2_valid, add_31_in1_valid}), .ready_in_bus({add_31_in2_ready, add_31_in1_ready}), 
		.data_out_bus({add_31_out1_data}), .valid_out_bus({add_31_out1_valid}), .ready_out_bus({add_31_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) const_node_cst_10
		(.clk(cst_10_clk), .rst(cst_10_rst),
		.data_in_bus({4'd8}), .valid_in_bus({cst_10_in1_valid}), .ready_in_bus({cst_10_in1_ready}), 
		.data_out_bus({cst_10_out1_data}), .valid_out_bus({cst_10_out1_valid}), .ready_out_bus({cst_10_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_32
		(.clk(icmp_32_clk), .rst(icmp_32_rst),
		.data_in_bus({icmp_32_in2_data, icmp_32_in1_data}), .valid_in_bus({icmp_32_in2_valid, icmp_32_in1_valid}), .ready_in_bus({icmp_32_in2_ready, icmp_32_in1_ready}), 
		.data_out_bus({icmp_32_out1_data}), .valid_out_bus({icmp_32_out1_valid}), .ready_out_bus({icmp_32_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n5
		(.clk(phi_n5_clk), .rst(phi_n5_rst),
		.data_in_bus({phi_n5_in1_data}), .valid_in_bus({phi_n5_in1_valid}), .ready_in_bus({phi_n5_in1_ready}), 
		.data_out_bus({phi_n5_out1_data}), .valid_out_bus({phi_n5_out1_valid}), .ready_out_bus({phi_n5_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n6
		(.clk(phi_n6_clk), .rst(phi_n6_rst),
		.data_in_bus({phi_n6_in1_data}), .valid_in_bus({phi_n6_in1_valid}), .ready_in_bus({phi_n6_in1_ready}), 
		.data_out_bus({phi_n6_out1_data}), .valid_out_bus({phi_n6_out1_valid}), .ready_out_bus({phi_n6_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n7
		(.clk(phi_n7_clk), .rst(phi_n7_rst),
		.data_in_bus({phi_n7_in1_data}), .valid_in_bus({phi_n7_in1_valid}), .ready_in_bus({phi_n7_in1_ready}), 
		.data_out_bus({phi_n7_out1_data}), .valid_out_bus({phi_n7_out1_valid}), .ready_out_bus({phi_n7_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_4
		(.clk(fork_4_clk), .rst(fork_4_rst),
		.data_in_bus({fork_4_in1_data}), .valid_in_bus({fork_4_in1_valid}), .ready_in_bus({fork_4_in1_ready}), 
		.data_out_bus({fork_4_out2_data, fork_4_out1_data}), .valid_out_bus({fork_4_out2_valid, fork_4_out1_valid}), .ready_out_bus({fork_4_out2_ready, fork_4_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_21
		(.clk(fork_21_clk), .rst(fork_21_rst),
		.data_in_bus({fork_21_in1_data}), .valid_in_bus({fork_21_in1_valid}), .ready_in_bus({fork_21_in1_ready}), 
		.data_out_bus({fork_21_out2_data, fork_21_out1_data}), .valid_out_bus({fork_21_out2_valid, fork_21_out1_valid}), .ready_out_bus({fork_21_out2_ready, fork_21_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_22
		(.clk(fork_22_clk), .rst(fork_22_rst),
		.data_in_bus({fork_22_in1_data}), .valid_in_bus({fork_22_in1_valid}), .ready_in_bus({fork_22_in1_ready}), 
		.data_out_bus({fork_22_out2_data, fork_22_out1_data}), .valid_out_bus({fork_22_out2_valid, fork_22_out1_valid}), .ready_out_bus({fork_22_out2_ready, fork_22_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_11
		(.clk(branch_11_clk), .rst(branch_11_rst),
		.data_in_bus({{3'b0, branch_11_in2_data}, branch_11_in1_data}), .valid_in_bus({branch_11_in2_valid, branch_11_in1_valid}), .ready_in_bus({branch_11_in2_ready, branch_11_in1_ready}), 
		.data_out_bus({branch_11_out2_data, branch_11_out1_data}), .valid_out_bus({branch_11_out2_valid, branch_11_out1_valid}), .ready_out_bus({branch_11_out2_ready, branch_11_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_12
		(.clk(branch_12_clk), .rst(branch_12_rst),
		.data_in_bus({{3'b0, branch_12_in2_data}, branch_12_in1_data}), .valid_in_bus({branch_12_in2_valid, branch_12_in1_valid}), .ready_in_bus({branch_12_in2_ready, branch_12_in1_ready}), 
		.data_out_bus({branch_12_out2_data, branch_12_out1_data}), .valid_out_bus({branch_12_out2_valid, branch_12_out1_valid}), .ready_out_bus({branch_12_out2_ready, branch_12_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_37
		(.clk(fork_37_clk), .rst(fork_37_rst),
		.data_in_bus({fork_37_in1_data}), .valid_in_bus({fork_37_in1_valid}), .ready_in_bus({fork_37_in1_ready}), 
		.data_out_bus({fork_37_out3_data, fork_37_out2_data, fork_37_out1_data}), .valid_out_bus({fork_37_out3_valid, fork_37_out2_valid, fork_37_out1_valid}), .ready_out_bus({fork_37_out3_ready, fork_37_out2_ready, fork_37_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_39
		(.clk(cst_39_clk), .rst(cst_39_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_39_in1_valid}), .ready_in_bus({cst_39_in1_ready}), 
		.data_out_bus({cst_39_out1_data}), .valid_out_bus({cst_39_out1_valid}), .ready_out_bus({cst_39_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_24
		(.clk(phiC_24_clk), .rst(phiC_24_rst),
		.data_in_bus({phiC_24_in1_data}), .valid_in_bus({phiC_24_in1_valid}), .ready_in_bus({phiC_24_in1_ready}), 
		.data_out_bus({phiC_24_out1_data}), .valid_out_bus({phiC_24_out1_valid}), .ready_out_bus({phiC_24_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_57
		(.clk(forkC_57_clk), .rst(forkC_57_rst),
		.data_in_bus({forkC_57_in1_data}), .valid_in_bus({forkC_57_in1_valid}), .ready_in_bus({forkC_57_in1_ready}), 
		.data_out_bus({forkC_57_out2_data, forkC_57_out1_data}), .valid_out_bus({forkC_57_out2_valid, forkC_57_out1_valid}), .ready_out_bus({forkC_57_out2_ready, forkC_57_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_46
		(.clk(branchC_46_clk), .rst(branchC_46_rst),
		.data_in_bus({{branchC_46_in2_data}, branchC_46_in1_data}), .valid_in_bus({branchC_46_in2_valid, branchC_46_in1_valid}), .ready_in_bus({branchC_46_in2_ready, branchC_46_in1_ready}), 
		.data_out_bus({branchC_46_out2_data, branchC_46_out1_data}), .valid_out_bus({branchC_46_out2_valid, branchC_46_out1_valid}), .ready_out_bus({branchC_46_out2_ready, branchC_46_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_5
		(.clk(source_5_clk), .rst(source_5_rst),
		.data_out_bus({source_5_out1_data}), .valid_out_bus({source_5_out1_valid}), .ready_out_bus({source_5_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_6
		(.clk(source_6_clk), .rst(source_6_rst),
		.data_out_bus({source_6_out1_data}), .valid_out_bus({source_6_out1_valid}), .ready_out_bus({source_6_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(4))source_node_source_7
		(.clk(source_7_clk), .rst(source_7_rst),
		.data_out_bus({source_7_out1_data}), .valid_out_bus({source_7_out1_valid}), .ready_out_bus({source_7_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block1
		(.clk(brCst_block1_clk), .rst(brCst_block1_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block1_in1_valid}), .ready_in_bus({brCst_block1_in1_ready}), 
		.data_out_bus({brCst_block1_out1_data}), .valid_out_bus({brCst_block1_out1_valid}), .ready_out_bus({brCst_block1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_0
		(.clk(cst_0_clk), .rst(cst_0_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_0_in1_valid}), .ready_in_bus({cst_0_in1_ready}), 
		.data_out_bus({cst_0_out1_data}), .valid_out_bus({cst_0_out1_valid}), .ready_out_bus({cst_0_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_0
		(.clk(branch_0_clk), .rst(branch_0_rst),
		.data_in_bus({{branch_0_in2_data}, branch_0_in1_data}), .valid_in_bus({branch_0_in2_valid, branch_0_in1_valid}), .ready_in_bus({branch_0_in2_ready, branch_0_in1_ready}), 
		.data_out_bus({branch_0_out2_data, branch_0_out1_data}), .valid_out_bus({branch_0_out2_valid, branch_0_out1_valid}), .ready_out_bus({branch_0_out2_ready, branch_0_out1_ready}));

	start_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) start_node_start_0
		(.clk(start_0_clk), .rst(start_0_rst),
		.data_in_bus({start_0_in1_data}), .valid_in_bus({start_0_in1_valid}), .ready_in_bus({start_0_in1_ready}), 
		.data_out_bus({start_0_out1_data}), .valid_out_bus({start_0_out1_valid}), .ready_out_bus({start_0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_52
		(.clk(forkC_52_clk), .rst(forkC_52_rst),
		.data_in_bus({forkC_52_in1_data}), .valid_in_bus({forkC_52_in1_valid}), .ready_in_bus({forkC_52_in1_ready}), 
		.data_out_bus({forkC_52_out3_data, forkC_52_out2_data, forkC_52_out1_data}), .valid_out_bus({forkC_52_out3_valid, forkC_52_out2_valid, forkC_52_out1_valid}), .ready_out_bus({forkC_52_out3_ready, forkC_52_out2_ready, forkC_52_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_42
		(.clk(branchC_42_clk), .rst(branchC_42_rst),
		.data_in_bus({{branchC_42_in2_data}, branchC_42_in1_data}), .valid_in_bus({branchC_42_in2_valid, branchC_42_in1_valid}), .ready_in_bus({branchC_42_in2_ready, branchC_42_in1_ready}), 
		.data_out_bus({branchC_42_out2_data, branchC_42_out1_data}), .valid_out_bus({branchC_42_out2_valid, branchC_42_out1_valid}), .ready_out_bus({branchC_42_out2_ready, branchC_42_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_53
		(.clk(fork_53_clk), .rst(fork_53_rst),
		.data_in_bus({fork_53_in1_data}), .valid_in_bus({fork_53_in1_valid}), .ready_in_bus({fork_53_in1_ready}), 
		.data_out_bus({fork_53_out2_data, fork_53_out1_data}), .valid_out_bus({fork_53_out2_valid, fork_53_out1_valid}), .ready_out_bus({fork_53_out2_ready, fork_53_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4), .COND_SIZE(1)) mux_node_phi_77
		(.clk(phi_77_clk), .rst(phi_77_rst),
		.data_in_bus({{3'b0, phi_77_in1_data}, phi_77_in3_data, phi_77_in2_data}), .valid_in_bus({phi_77_in1_valid, phi_77_in3_valid, phi_77_in2_valid}), .ready_in_bus({phi_77_in1_ready, phi_77_in3_ready, phi_77_in2_ready}), 
		.data_out_bus({phi_77_out1_data}), .valid_out_bus({phi_77_out1_valid}), .ready_out_bus({phi_77_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_28
		(.clk(cst_28_clk), .rst(cst_28_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_28_in1_valid}), .ready_in_bus({cst_28_in1_ready}), 
		.data_out_bus({cst_28_out1_data}), .valid_out_bus({cst_28_out1_valid}), .ready_out_bus({cst_28_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_78
		(.clk(shl_78_clk), .rst(shl_78_rst),
		.data_in_bus({shl_78_in2_data, shl_78_in1_data}), .valid_in_bus({shl_78_in2_valid, shl_78_in1_valid}), .ready_in_bus({shl_78_in2_ready, shl_78_in1_ready}), 
		.data_out_bus({shl_78_out1_data}), .valid_out_bus({shl_78_out1_valid}), .ready_out_bus({shl_78_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_79
		(.clk(add_79_clk), .rst(add_79_rst),
		.data_in_bus({add_79_in2_data, add_79_in1_data}), .valid_in_bus({add_79_in2_valid, add_79_in1_valid}), .ready_in_bus({add_79_in2_ready, add_79_in1_ready}), 
		.data_out_bus({add_79_out1_data}), .valid_out_bus({add_79_out1_valid}), .ready_out_bus({add_79_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_load_op_load_82
		(.clk(load_82_clk), .rst(load_82_rst),
		.data_in_bus({load_82_in1_data}), .address_in_bus({load_82_in2_data}), .valid_in_bus({load_82_in2_valid, load_82_in1_valid}), .ready_in_bus({load_82_in2_ready, load_82_in1_ready}), 
		.data_out_bus({load_82_out1_data}), .address_out_bus({load_82_out2_data}), .valid_out_bus({load_82_out2_valid, load_82_out1_valid}), .ready_out_bus({load_82_out2_ready, load_82_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block15
		(.clk(brCst_block15_clk), .rst(brCst_block15_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block15_in1_valid}), .ready_in_bus({brCst_block15_in1_ready}), 
		.data_out_bus({brCst_block15_out1_data}), .valid_out_bus({brCst_block15_out1_valid}), .ready_out_bus({brCst_block15_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_29
		(.clk(cst_29_clk), .rst(cst_29_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_29_in1_valid}), .ready_in_bus({cst_29_in1_ready}), 
		.data_out_bus({cst_29_out1_data}), .valid_out_bus({cst_29_out1_valid}), .ready_out_bus({cst_29_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n15
		(.clk(phi_n15_clk), .rst(phi_n15_rst),
		.data_in_bus({phi_n15_in2_data, phi_n15_in1_data}), .valid_in_bus({phi_n15_in2_valid, phi_n15_in1_valid}), .ready_in_bus({phi_n15_in2_ready, phi_n15_in1_ready}), 
		.data_out_bus({phi_n15_out1_data}), .valid_out_bus({phi_n15_out1_valid}), .ready_out_bus({phi_n15_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_12
		(.clk(fork_12_clk), .rst(fork_12_rst),
		.data_in_bus({fork_12_in1_data}), .valid_in_bus({fork_12_in1_valid}), .ready_in_bus({fork_12_in1_ready}), 
		.data_out_bus({fork_12_out2_data, fork_12_out1_data}), .valid_out_bus({fork_12_out2_valid, fork_12_out1_valid}), .ready_out_bus({fork_12_out2_ready, fork_12_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_28
		(.clk(fork_28_clk), .rst(fork_28_rst),
		.data_in_bus({fork_28_in1_data}), .valid_in_bus({fork_28_in1_valid}), .ready_in_bus({fork_28_in1_ready}), 
		.data_out_bus({fork_28_out2_data, fork_28_out1_data}), .valid_out_bus({fork_28_out2_valid, fork_28_out1_valid}), .ready_out_bus({fork_28_out2_ready, fork_28_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_31
		(.clk(branch_31_clk), .rst(branch_31_rst),
		.data_in_bus({{31'b0, branch_31_in2_data}, branch_31_in1_data}), .valid_in_bus({branch_31_in2_valid, branch_31_in1_valid}), .ready_in_bus({branch_31_in2_ready, branch_31_in1_ready}), 
		.data_out_bus({branch_31_out2_data, branch_31_out1_data}), .valid_out_bus({branch_31_out2_valid, branch_31_out1_valid}), .ready_out_bus({branch_31_out2_ready, branch_31_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_32
		(.clk(branch_32_clk), .rst(branch_32_rst),
		.data_in_bus({{branch_32_in2_data}, branch_32_in1_data}), .valid_in_bus({branch_32_in2_valid, branch_32_in1_valid}), .ready_in_bus({branch_32_in2_ready, branch_32_in1_ready}), 
		.data_out_bus({branch_32_out2_data, branch_32_out1_data}), .valid_out_bus({branch_32_out2_valid, branch_32_out1_valid}), .ready_out_bus({branch_32_out2_ready, branch_32_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_33
		(.clk(branch_33_clk), .rst(branch_33_rst),
		.data_in_bus({{3'b0, branch_33_in2_data}, branch_33_in1_data}), .valid_in_bus({branch_33_in2_valid, branch_33_in1_valid}), .ready_in_bus({branch_33_in2_ready, branch_33_in1_ready}), 
		.data_out_bus({branch_33_out2_data, branch_33_out1_data}), .valid_out_bus({branch_33_out2_valid, branch_33_out1_valid}), .ready_out_bus({branch_33_out2_ready, branch_33_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_34
		(.clk(branch_34_clk), .rst(branch_34_rst),
		.data_in_bus({{3'b0, branch_34_in2_data}, branch_34_in1_data}), .valid_in_bus({branch_34_in2_valid, branch_34_in1_valid}), .ready_in_bus({branch_34_in2_ready, branch_34_in1_ready}), 
		.data_out_bus({branch_34_out2_data, branch_34_out1_data}), .valid_out_bus({branch_34_out2_valid, branch_34_out1_valid}), .ready_out_bus({branch_34_out2_ready, branch_34_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_47
		(.clk(fork_47_clk), .rst(fork_47_rst),
		.data_in_bus({fork_47_in1_data}), .valid_in_bus({fork_47_in1_valid}), .ready_in_bus({fork_47_in1_ready}), 
		.data_out_bus({fork_47_out5_data, fork_47_out4_data, fork_47_out3_data, fork_47_out2_data, fork_47_out1_data}), .valid_out_bus({fork_47_out5_valid, fork_47_out4_valid, fork_47_out3_valid, fork_47_out2_valid, fork_47_out1_valid}), .ready_out_bus({fork_47_out5_ready, fork_47_out4_ready, fork_47_out3_ready, fork_47_out2_ready, fork_47_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_34
		(.clk(phiC_34_clk), .rst(phiC_34_rst),
		.data_in_bus({phiC_34_in2_data, phiC_34_in1_data}), .valid_in_bus({phiC_34_in2_valid, phiC_34_in1_valid}), .ready_in_bus({phiC_34_in2_ready, phiC_34_in1_ready}), 
		.data_out_bus({phiC_34_out2_data, phiC_34_out1_data}), .valid_out_bus({phiC_34_out2_valid, phiC_34_out1_valid}), .ready_out_bus({phiC_34_out2_ready, phiC_34_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_71
		(.clk(forkC_71_clk), .rst(forkC_71_rst),
		.data_in_bus({forkC_71_in1_data}), .valid_in_bus({forkC_71_in1_valid}), .ready_in_bus({forkC_71_in1_ready}), 
		.data_out_bus({forkC_71_out3_data, forkC_71_out2_data, forkC_71_out1_data}), .valid_out_bus({forkC_71_out3_valid, forkC_71_out2_valid, forkC_71_out1_valid}), .ready_out_bus({forkC_71_out3_ready, forkC_71_out2_ready, forkC_71_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_56
		(.clk(branchC_56_clk), .rst(branchC_56_rst),
		.data_in_bus({{branchC_56_in2_data}, branchC_56_in1_data}), .valid_in_bus({branchC_56_in2_valid, branchC_56_in1_valid}), .ready_in_bus({branchC_56_in2_ready, branchC_56_in1_ready}), 
		.data_out_bus({branchC_56_out2_data, branchC_56_out1_data}), .valid_out_bus({branchC_56_out2_valid, branchC_56_out1_valid}), .ready_out_bus({branchC_56_out2_ready, branchC_56_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_20
		(.clk(source_20_clk), .rst(source_20_rst),
		.data_out_bus({source_20_out1_data}), .valid_out_bus({source_20_out1_valid}), .ready_out_bus({source_20_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4), .COND_SIZE(1)) mux_node_phi_38
		(.clk(phi_38_clk), .rst(phi_38_rst),
		.data_in_bus({{3'b0, phi_38_in1_data}, phi_38_in3_data, phi_38_in2_data}), .valid_in_bus({phi_38_in1_valid, phi_38_in3_valid, phi_38_in2_valid}), .ready_in_bus({phi_38_in1_ready, phi_38_in3_ready, phi_38_in2_ready}), 
		.data_out_bus({phi_38_out1_data}), .valid_out_bus({phi_38_out1_valid}), .ready_out_bus({phi_38_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block8
		(.clk(brCst_block8_clk), .rst(brCst_block8_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block8_in1_valid}), .ready_in_bus({brCst_block8_in1_ready}), 
		.data_out_bus({brCst_block8_out1_data}), .valid_out_bus({brCst_block8_out1_valid}), .ready_out_bus({brCst_block8_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_14
		(.clk(cst_14_clk), .rst(cst_14_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_14_in1_valid}), .ready_in_bus({cst_14_in1_ready}), 
		.data_out_bus({cst_14_out1_data}), .valid_out_bus({cst_14_out1_valid}), .ready_out_bus({cst_14_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_15
		(.clk(branch_15_clk), .rst(branch_15_rst),
		.data_in_bus({{branch_15_in2_data}, branch_15_in1_data}), .valid_in_bus({branch_15_in2_valid, branch_15_in1_valid}), .ready_in_bus({branch_15_in2_ready, branch_15_in1_ready}), 
		.data_out_bus({branch_15_out2_data, branch_15_out1_data}), .valid_out_bus({branch_15_out2_valid, branch_15_out1_valid}), .ready_out_bus({branch_15_out2_ready, branch_15_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_16
		(.clk(branch_16_clk), .rst(branch_16_rst),
		.data_in_bus({{3'b0, branch_16_in2_data}, branch_16_in1_data}), .valid_in_bus({branch_16_in2_valid, branch_16_in1_valid}), .ready_in_bus({branch_16_in2_ready, branch_16_in1_ready}), 
		.data_out_bus({branch_16_out2_data, branch_16_out1_data}), .valid_out_bus({branch_16_out2_valid, branch_16_out1_valid}), .ready_out_bus({branch_16_out2_ready, branch_16_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_40
		(.clk(fork_40_clk), .rst(fork_40_rst),
		.data_in_bus({fork_40_in1_data}), .valid_in_bus({fork_40_in1_valid}), .ready_in_bus({fork_40_in1_ready}), 
		.data_out_bus({fork_40_out3_data, fork_40_out2_data, fork_40_out1_data}), .valid_out_bus({fork_40_out3_valid, fork_40_out2_valid, fork_40_out1_valid}), .ready_out_bus({fork_40_out3_ready, fork_40_out2_ready, fork_40_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_27
		(.clk(phiC_27_clk), .rst(phiC_27_rst),
		.data_in_bus({phiC_27_in2_data, phiC_27_in1_data}), .valid_in_bus({phiC_27_in2_valid, phiC_27_in1_valid}), .ready_in_bus({phiC_27_in2_ready, phiC_27_in1_ready}), 
		.data_out_bus({phiC_27_out2_data, phiC_27_out1_data}), .valid_out_bus({phiC_27_out2_valid, phiC_27_out1_valid}), .ready_out_bus({phiC_27_out2_ready, phiC_27_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_62
		(.clk(forkC_62_clk), .rst(forkC_62_rst),
		.data_in_bus({forkC_62_in1_data}), .valid_in_bus({forkC_62_in1_valid}), .ready_in_bus({forkC_62_in1_ready}), 
		.data_out_bus({forkC_62_out3_data, forkC_62_out2_data, forkC_62_out1_data}), .valid_out_bus({forkC_62_out3_valid, forkC_62_out2_valid, forkC_62_out1_valid}), .ready_out_bus({forkC_62_out3_ready, forkC_62_out2_ready, forkC_62_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_49
		(.clk(branchC_49_clk), .rst(branchC_49_rst),
		.data_in_bus({{branchC_49_in2_data}, branchC_49_in1_data}), .valid_in_bus({branchC_49_in2_valid, branchC_49_in1_valid}), .ready_in_bus({branchC_49_in2_ready, branchC_49_in1_ready}), 
		.data_out_bus({branchC_49_out2_data, branchC_49_out1_data}), .valid_out_bus({branchC_49_out2_valid, branchC_49_out1_valid}), .ready_out_bus({branchC_49_out2_ready, branchC_49_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_11
		(.clk(cst_11_clk), .rst(cst_11_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_11_in1_valid}), .ready_in_bus({cst_11_in1_ready}), 
		.data_out_bus({cst_11_out1_data}), .valid_out_bus({cst_11_out1_valid}), .ready_out_bus({cst_11_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) add_op_add_34
		(.clk(add_34_clk), .rst(add_34_rst),
		.data_in_bus({add_34_in2_data, add_34_in1_data}), .valid_in_bus({add_34_in2_valid, add_34_in1_valid}), .ready_in_bus({add_34_in2_ready, add_34_in1_ready}), 
		.data_out_bus({add_34_out1_data}), .valid_out_bus({add_34_out1_valid}), .ready_out_bus({add_34_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) const_node_cst_12
		(.clk(cst_12_clk), .rst(cst_12_rst),
		.data_in_bus({4'd8}), .valid_in_bus({cst_12_in1_valid}), .ready_in_bus({cst_12_in1_ready}), 
		.data_out_bus({cst_12_out1_data}), .valid_out_bus({cst_12_out1_valid}), .ready_out_bus({cst_12_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_35
		(.clk(icmp_35_clk), .rst(icmp_35_rst),
		.data_in_bus({icmp_35_in2_data, icmp_35_in1_data}), .valid_in_bus({icmp_35_in2_valid, icmp_35_in1_valid}), .ready_in_bus({icmp_35_in2_ready, icmp_35_in1_ready}), 
		.data_out_bus({icmp_35_out1_data}), .valid_out_bus({icmp_35_out1_valid}), .ready_out_bus({icmp_35_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n3
		(.clk(phi_n3_clk), .rst(phi_n3_rst),
		.data_in_bus({phi_n3_in1_data}), .valid_in_bus({phi_n3_in1_valid}), .ready_in_bus({phi_n3_in1_ready}), 
		.data_out_bus({phi_n3_out1_data}), .valid_out_bus({phi_n3_out1_valid}), .ready_out_bus({phi_n3_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_5
		(.clk(fork_5_clk), .rst(fork_5_rst),
		.data_in_bus({fork_5_in1_data}), .valid_in_bus({fork_5_in1_valid}), .ready_in_bus({fork_5_in1_ready}), 
		.data_out_bus({fork_5_out2_data, fork_5_out1_data}), .valid_out_bus({fork_5_out2_valid, fork_5_out1_valid}), .ready_out_bus({fork_5_out2_ready, fork_5_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_13
		(.clk(branch_13_clk), .rst(branch_13_rst),
		.data_in_bus({{3'b0, branch_13_in2_data}, branch_13_in1_data}), .valid_in_bus({branch_13_in2_valid, branch_13_in1_valid}), .ready_in_bus({branch_13_in2_ready, branch_13_in1_ready}), 
		.data_out_bus({branch_13_out2_data, branch_13_out1_data}), .valid_out_bus({branch_13_out2_valid, branch_13_out1_valid}), .ready_out_bus({branch_13_out2_ready, branch_13_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_25
		(.clk(phiC_25_clk), .rst(phiC_25_rst),
		.data_in_bus({phiC_25_in1_data}), .valid_in_bus({phiC_25_in1_valid}), .ready_in_bus({phiC_25_in1_ready}), 
		.data_out_bus({phiC_25_out1_data}), .valid_out_bus({phiC_25_out1_valid}), .ready_out_bus({phiC_25_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_47
		(.clk(branchC_47_clk), .rst(branchC_47_rst),
		.data_in_bus({{branchC_47_in2_data}, branchC_47_in1_data}), .valid_in_bus({branchC_47_in2_valid, branchC_47_in1_valid}), .ready_in_bus({branchC_47_in2_ready, branchC_47_in1_ready}), 
		.data_out_bus({branchC_47_out2_data, branchC_47_out1_data}), .valid_out_bus({branchC_47_out2_valid, branchC_47_out1_valid}), .ready_out_bus({branchC_47_out2_ready, branchC_47_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_59
		(.clk(fork_59_clk), .rst(fork_59_rst),
		.data_in_bus({fork_59_in1_data}), .valid_in_bus({fork_59_in1_valid}), .ready_in_bus({fork_59_in1_ready}), 
		.data_out_bus({fork_59_out2_data, fork_59_out1_data}), .valid_out_bus({fork_59_out2_valid, fork_59_out1_valid}), .ready_out_bus({fork_59_out2_ready, fork_59_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_8
		(.clk(source_8_clk), .rst(source_8_rst),
		.data_out_bus({source_8_out1_data}), .valid_out_bus({source_8_out1_valid}), .ready_out_bus({source_8_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(4))source_node_source_9
		(.clk(source_9_clk), .rst(source_9_rst),
		.data_out_bus({source_9_out1_data}), .valid_out_bus({source_9_out1_valid}), .ready_out_bus({source_9_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_34
		(.clk(cst_34_clk), .rst(cst_34_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_34_in1_valid}), .ready_in_bus({cst_34_in1_ready}), 
		.data_out_bus({cst_34_out1_data}), .valid_out_bus({cst_34_out1_valid}), .ready_out_bus({cst_34_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_101
		(.clk(shl_101_clk), .rst(shl_101_rst),
		.data_in_bus({shl_101_in2_data, shl_101_in1_data}), .valid_in_bus({shl_101_in2_valid, shl_101_in1_valid}), .ready_in_bus({shl_101_in2_ready, shl_101_in1_ready}), 
		.data_out_bus({shl_101_out1_data}), .valid_out_bus({shl_101_out1_valid}), .ready_out_bus({shl_101_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_102
		(.clk(add_102_clk), .rst(add_102_rst),
		.data_in_bus({add_102_in2_data, add_102_in1_data}), .valid_in_bus({add_102_in2_valid, add_102_in1_valid}), .ready_in_bus({add_102_in2_ready, add_102_in1_ready}), 
		.data_out_bus({add_102_out1_data}), .valid_out_bus({add_102_out1_valid}), .ready_out_bus({add_102_out1_ready}));

	mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_store_op_store_2
		(.clk(store_2_clk), .rst(store_2_rst),
		.data_in_bus({store_2_in1_data}), .address_in_bus({store_2_in2_data}), .valid_in_bus({store_2_in2_valid, store_2_in1_valid}), .ready_in_bus({store_2_in2_ready, store_2_in1_ready}), 
		.data_out_bus({store_2_out1_data}), .address_out_bus({store_2_out2_data}), .valid_out_bus({store_2_out2_valid, store_2_out1_valid}), .ready_out_bus({store_2_out2_ready, store_2_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_35
		(.clk(cst_35_clk), .rst(cst_35_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_35_in1_valid}), .ready_in_bus({cst_35_in1_ready}), 
		.data_out_bus({cst_35_out1_data}), .valid_out_bus({cst_35_out1_valid}), .ready_out_bus({cst_35_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) add_op_add_105
		(.clk(add_105_clk), .rst(add_105_rst),
		.data_in_bus({add_105_in2_data, add_105_in1_data}), .valid_in_bus({add_105_in2_valid, add_105_in1_valid}), .ready_in_bus({add_105_in2_ready, add_105_in1_ready}), 
		.data_out_bus({add_105_out1_data}), .valid_out_bus({add_105_out1_valid}), .ready_out_bus({add_105_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) const_node_cst_36
		(.clk(cst_36_clk), .rst(cst_36_rst),
		.data_in_bus({4'd8}), .valid_in_bus({cst_36_in1_valid}), .ready_in_bus({cst_36_in1_ready}), 
		.data_out_bus({cst_36_out1_data}), .valid_out_bus({cst_36_out1_valid}), .ready_out_bus({cst_36_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_106
		(.clk(icmp_106_clk), .rst(icmp_106_rst),
		.data_in_bus({icmp_106_in2_data, icmp_106_in1_data}), .valid_in_bus({icmp_106_in2_valid, icmp_106_in1_valid}), .ready_in_bus({icmp_106_in2_ready, icmp_106_in1_ready}), 
		.data_out_bus({icmp_106_out1_data}), .valid_out_bus({icmp_106_out1_valid}), .ready_out_bus({icmp_106_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n16
		(.clk(phi_n16_clk), .rst(phi_n16_rst),
		.data_in_bus({phi_n16_in1_data}), .valid_in_bus({phi_n16_in1_valid}), .ready_in_bus({phi_n16_in1_ready}), 
		.data_out_bus({phi_n16_out1_data}), .valid_out_bus({phi_n16_out1_valid}), .ready_out_bus({phi_n16_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n17
		(.clk(phi_n17_clk), .rst(phi_n17_rst),
		.data_in_bus({phi_n17_in1_data}), .valid_in_bus({phi_n17_in1_valid}), .ready_in_bus({phi_n17_in1_ready}), 
		.data_out_bus({phi_n17_out1_data}), .valid_out_bus({phi_n17_out1_valid}), .ready_out_bus({phi_n17_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n18
		(.clk(phi_n18_clk), .rst(phi_n18_rst),
		.data_in_bus({phi_n18_in1_data}), .valid_in_bus({phi_n18_in1_valid}), .ready_in_bus({phi_n18_in1_ready}), 
		.data_out_bus({phi_n18_out1_data}), .valid_out_bus({phi_n18_out1_valid}), .ready_out_bus({phi_n18_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_16
		(.clk(fork_16_clk), .rst(fork_16_rst),
		.data_in_bus({fork_16_in1_data}), .valid_in_bus({fork_16_in1_valid}), .ready_in_bus({fork_16_in1_ready}), 
		.data_out_bus({fork_16_out2_data, fork_16_out1_data}), .valid_out_bus({fork_16_out2_valid, fork_16_out1_valid}), .ready_out_bus({fork_16_out2_ready, fork_16_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_29
		(.clk(fork_29_clk), .rst(fork_29_rst),
		.data_in_bus({fork_29_in1_data}), .valid_in_bus({fork_29_in1_valid}), .ready_in_bus({fork_29_in1_ready}), 
		.data_out_bus({fork_29_out2_data, fork_29_out1_data}), .valid_out_bus({fork_29_out2_valid, fork_29_out1_valid}), .ready_out_bus({fork_29_out2_ready, fork_29_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_30
		(.clk(fork_30_clk), .rst(fork_30_rst),
		.data_in_bus({fork_30_in1_data}), .valid_in_bus({fork_30_in1_valid}), .ready_in_bus({fork_30_in1_ready}), 
		.data_out_bus({fork_30_out2_data, fork_30_out1_data}), .valid_out_bus({fork_30_out2_valid, fork_30_out1_valid}), .ready_out_bus({fork_30_out2_ready, fork_30_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_39
		(.clk(branch_39_clk), .rst(branch_39_rst),
		.data_in_bus({{3'b0, branch_39_in2_data}, branch_39_in1_data}), .valid_in_bus({branch_39_in2_valid, branch_39_in1_valid}), .ready_in_bus({branch_39_in2_ready, branch_39_in1_ready}), 
		.data_out_bus({branch_39_out2_data, branch_39_out1_data}), .valid_out_bus({branch_39_out2_valid, branch_39_out1_valid}), .ready_out_bus({branch_39_out2_ready, branch_39_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_40
		(.clk(branch_40_clk), .rst(branch_40_rst),
		.data_in_bus({{3'b0, branch_40_in2_data}, branch_40_in1_data}), .valid_in_bus({branch_40_in2_valid, branch_40_in1_valid}), .ready_in_bus({branch_40_in2_ready, branch_40_in1_ready}), 
		.data_out_bus({branch_40_out2_data, branch_40_out1_data}), .valid_out_bus({branch_40_out2_valid, branch_40_out1_valid}), .ready_out_bus({branch_40_out2_ready, branch_40_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_49
		(.clk(fork_49_clk), .rst(fork_49_rst),
		.data_in_bus({fork_49_in1_data}), .valid_in_bus({fork_49_in1_valid}), .ready_in_bus({fork_49_in1_ready}), 
		.data_out_bus({fork_49_out3_data, fork_49_out2_data, fork_49_out1_data}), .valid_out_bus({fork_49_out3_valid, fork_49_out2_valid, fork_49_out1_valid}), .ready_out_bus({fork_49_out3_ready, fork_49_out2_ready, fork_49_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_41
		(.clk(cst_41_clk), .rst(cst_41_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_41_in1_valid}), .ready_in_bus({cst_41_in1_ready}), 
		.data_out_bus({cst_41_out1_data}), .valid_out_bus({cst_41_out1_valid}), .ready_out_bus({cst_41_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_36
		(.clk(phiC_36_clk), .rst(phiC_36_rst),
		.data_in_bus({phiC_36_in1_data}), .valid_in_bus({phiC_36_in1_valid}), .ready_in_bus({phiC_36_in1_ready}), 
		.data_out_bus({phiC_36_out1_data}), .valid_out_bus({phiC_36_out1_valid}), .ready_out_bus({phiC_36_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_73
		(.clk(forkC_73_clk), .rst(forkC_73_rst),
		.data_in_bus({forkC_73_in1_data}), .valid_in_bus({forkC_73_in1_valid}), .ready_in_bus({forkC_73_in1_ready}), 
		.data_out_bus({forkC_73_out2_data, forkC_73_out1_data}), .valid_out_bus({forkC_73_out2_valid, forkC_73_out1_valid}), .ready_out_bus({forkC_73_out2_ready, forkC_73_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_58
		(.clk(branchC_58_clk), .rst(branchC_58_rst),
		.data_in_bus({{branchC_58_in2_data}, branchC_58_in1_data}), .valid_in_bus({branchC_58_in2_valid, branchC_58_in1_valid}), .ready_in_bus({branchC_58_in2_ready, branchC_58_in1_ready}), 
		.data_out_bus({branchC_58_out2_data, branchC_58_out1_data}), .valid_out_bus({branchC_58_out2_valid, branchC_58_out1_valid}), .ready_out_bus({branchC_58_out2_ready, branchC_58_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_25
		(.clk(source_25_clk), .rst(source_25_rst),
		.data_out_bus({source_25_out1_data}), .valid_out_bus({source_25_out1_valid}), .ready_out_bus({source_25_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_26
		(.clk(source_26_clk), .rst(source_26_rst),
		.data_out_bus({source_26_out1_data}), .valid_out_bus({source_26_out1_valid}), .ready_out_bus({source_26_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(4))source_node_source_27
		(.clk(source_27_clk), .rst(source_27_rst),
		.data_out_bus({source_27_out1_data}), .valid_out_bus({source_27_out1_valid}), .ready_out_bus({source_27_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_21
		(.clk(cst_21_clk), .rst(cst_21_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_21_in1_valid}), .ready_in_bus({cst_21_in1_ready}), 
		.data_out_bus({cst_21_out1_data}), .valid_out_bus({cst_21_out1_valid}), .ready_out_bus({cst_21_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_64
		(.clk(shl_64_clk), .rst(shl_64_rst),
		.data_in_bus({shl_64_in2_data, shl_64_in1_data}), .valid_in_bus({shl_64_in2_valid, shl_64_in1_valid}), .ready_in_bus({shl_64_in2_ready, shl_64_in1_ready}), 
		.data_out_bus({shl_64_out1_data}), .valid_out_bus({shl_64_out1_valid}), .ready_out_bus({shl_64_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_65
		(.clk(add_65_clk), .rst(add_65_rst),
		.data_in_bus({add_65_in2_data, add_65_in1_data}), .valid_in_bus({add_65_in2_valid, add_65_in1_valid}), .ready_in_bus({add_65_in2_ready, add_65_in1_ready}), 
		.data_out_bus({add_65_out1_data}), .valid_out_bus({add_65_out1_valid}), .ready_out_bus({add_65_out1_ready}));

	mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_store_op_store_1
		(.clk(store_1_clk), .rst(store_1_rst),
		.data_in_bus({store_1_in1_data}), .address_in_bus({store_1_in2_data}), .valid_in_bus({store_1_in2_valid, store_1_in1_valid}), .ready_in_bus({store_1_in2_ready, store_1_in1_ready}), 
		.data_out_bus({store_1_out1_data}), .address_out_bus({store_1_out2_data}), .valid_out_bus({store_1_out2_valid, store_1_out1_valid}), .ready_out_bus({store_1_out2_ready, store_1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_22
		(.clk(cst_22_clk), .rst(cst_22_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_22_in1_valid}), .ready_in_bus({cst_22_in1_ready}), 
		.data_out_bus({cst_22_out1_data}), .valid_out_bus({cst_22_out1_valid}), .ready_out_bus({cst_22_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) add_op_add_68
		(.clk(add_68_clk), .rst(add_68_rst),
		.data_in_bus({add_68_in2_data, add_68_in1_data}), .valid_in_bus({add_68_in2_valid, add_68_in1_valid}), .ready_in_bus({add_68_in2_ready, add_68_in1_ready}), 
		.data_out_bus({add_68_out1_data}), .valid_out_bus({add_68_out1_valid}), .ready_out_bus({add_68_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) const_node_cst_23
		(.clk(cst_23_clk), .rst(cst_23_rst),
		.data_in_bus({4'd8}), .valid_in_bus({cst_23_in1_valid}), .ready_in_bus({cst_23_in1_ready}), 
		.data_out_bus({cst_23_out1_data}), .valid_out_bus({cst_23_out1_valid}), .ready_out_bus({cst_23_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_69
		(.clk(icmp_69_clk), .rst(icmp_69_rst),
		.data_in_bus({icmp_69_in2_data, icmp_69_in1_data}), .valid_in_bus({icmp_69_in2_valid, icmp_69_in1_valid}), .ready_in_bus({icmp_69_in2_ready, icmp_69_in1_ready}), 
		.data_out_bus({icmp_69_out1_data}), .valid_out_bus({icmp_69_out1_valid}), .ready_out_bus({icmp_69_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n0
		(.clk(phi_n0_clk), .rst(phi_n0_rst),
		.data_in_bus({phi_n0_in1_data}), .valid_in_bus({phi_n0_in1_valid}), .ready_in_bus({phi_n0_in1_ready}), 
		.data_out_bus({phi_n0_out1_data}), .valid_out_bus({phi_n0_out1_valid}), .ready_out_bus({phi_n0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n1
		(.clk(phi_n1_clk), .rst(phi_n1_rst),
		.data_in_bus({phi_n1_in1_data}), .valid_in_bus({phi_n1_in1_valid}), .ready_in_bus({phi_n1_in1_ready}), 
		.data_out_bus({phi_n1_out1_data}), .valid_out_bus({phi_n1_out1_valid}), .ready_out_bus({phi_n1_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n2
		(.clk(phi_n2_clk), .rst(phi_n2_rst),
		.data_in_bus({phi_n2_in1_data}), .valid_in_bus({phi_n2_in1_valid}), .ready_in_bus({phi_n2_in1_ready}), 
		.data_out_bus({phi_n2_out1_data}), .valid_out_bus({phi_n2_out1_valid}), .ready_out_bus({phi_n2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_10
		(.clk(fork_10_clk), .rst(fork_10_rst),
		.data_in_bus({fork_10_in1_data}), .valid_in_bus({fork_10_in1_valid}), .ready_in_bus({fork_10_in1_ready}), 
		.data_out_bus({fork_10_out2_data, fork_10_out1_data}), .valid_out_bus({fork_10_out2_valid, fork_10_out1_valid}), .ready_out_bus({fork_10_out2_ready, fork_10_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_18
		(.clk(fork_18_clk), .rst(fork_18_rst),
		.data_in_bus({fork_18_in1_data}), .valid_in_bus({fork_18_in1_valid}), .ready_in_bus({fork_18_in1_ready}), 
		.data_out_bus({fork_18_out2_data, fork_18_out1_data}), .valid_out_bus({fork_18_out2_valid, fork_18_out1_valid}), .ready_out_bus({fork_18_out2_ready, fork_18_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_19
		(.clk(fork_19_clk), .rst(fork_19_rst),
		.data_in_bus({fork_19_in1_data}), .valid_in_bus({fork_19_in1_valid}), .ready_in_bus({fork_19_in1_ready}), 
		.data_out_bus({fork_19_out2_data, fork_19_out1_data}), .valid_out_bus({fork_19_out2_valid, fork_19_out1_valid}), .ready_out_bus({fork_19_out2_ready, fork_19_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_25
		(.clk(branch_25_clk), .rst(branch_25_rst),
		.data_in_bus({{3'b0, branch_25_in2_data}, branch_25_in1_data}), .valid_in_bus({branch_25_in2_valid, branch_25_in1_valid}), .ready_in_bus({branch_25_in2_ready, branch_25_in1_ready}), 
		.data_out_bus({branch_25_out2_data, branch_25_out1_data}), .valid_out_bus({branch_25_out2_valid, branch_25_out1_valid}), .ready_out_bus({branch_25_out2_ready, branch_25_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_26
		(.clk(branch_26_clk), .rst(branch_26_rst),
		.data_in_bus({{3'b0, branch_26_in2_data}, branch_26_in1_data}), .valid_in_bus({branch_26_in2_valid, branch_26_in1_valid}), .ready_in_bus({branch_26_in2_ready, branch_26_in1_ready}), 
		.data_out_bus({branch_26_out2_data, branch_26_out1_data}), .valid_out_bus({branch_26_out2_valid, branch_26_out1_valid}), .ready_out_bus({branch_26_out2_ready, branch_26_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_43
		(.clk(fork_43_clk), .rst(fork_43_rst),
		.data_in_bus({fork_43_in1_data}), .valid_in_bus({fork_43_in1_valid}), .ready_in_bus({fork_43_in1_ready}), 
		.data_out_bus({fork_43_out3_data, fork_43_out2_data, fork_43_out1_data}), .valid_out_bus({fork_43_out3_valid, fork_43_out2_valid, fork_43_out1_valid}), .ready_out_bus({fork_43_out3_ready, fork_43_out2_ready, fork_43_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_40
		(.clk(cst_40_clk), .rst(cst_40_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_40_in1_valid}), .ready_in_bus({cst_40_in1_ready}), 
		.data_out_bus({cst_40_out1_data}), .valid_out_bus({cst_40_out1_valid}), .ready_out_bus({cst_40_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_30
		(.clk(phiC_30_clk), .rst(phiC_30_rst),
		.data_in_bus({phiC_30_in1_data}), .valid_in_bus({phiC_30_in1_valid}), .ready_in_bus({phiC_30_in1_ready}), 
		.data_out_bus({phiC_30_out1_data}), .valid_out_bus({phiC_30_out1_valid}), .ready_out_bus({phiC_30_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_65
		(.clk(forkC_65_clk), .rst(forkC_65_rst),
		.data_in_bus({forkC_65_in1_data}), .valid_in_bus({forkC_65_in1_valid}), .ready_in_bus({forkC_65_in1_ready}), 
		.data_out_bus({forkC_65_out2_data, forkC_65_out1_data}), .valid_out_bus({forkC_65_out2_valid, forkC_65_out1_valid}), .ready_out_bus({forkC_65_out2_ready, forkC_65_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_52
		(.clk(branchC_52_clk), .rst(branchC_52_rst),
		.data_in_bus({{branchC_52_in2_data}, branchC_52_in1_data}), .valid_in_bus({branchC_52_in2_valid, branchC_52_in1_valid}), .ready_in_bus({branchC_52_in2_ready, branchC_52_in1_ready}), 
		.data_out_bus({branchC_52_out2_data, branchC_52_out1_data}), .valid_out_bus({branchC_52_out2_valid, branchC_52_out1_valid}), .ready_out_bus({branchC_52_out2_ready, branchC_52_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_15
		(.clk(source_15_clk), .rst(source_15_rst),
		.data_out_bus({source_15_out1_data}), .valid_out_bus({source_15_out1_valid}), .ready_out_bus({source_15_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_16
		(.clk(source_16_clk), .rst(source_16_rst),
		.data_out_bus({source_16_out1_data}), .valid_out_bus({source_16_out1_valid}), .ready_out_bus({source_16_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(4))source_node_source_17
		(.clk(source_17_clk), .rst(source_17_rst),
		.data_out_bus({source_17_out1_data}), .valid_out_bus({source_17_out1_valid}), .ready_out_bus({source_17_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4), .COND_SIZE(1)) mux_node_phi_40
		(.clk(phi_40_clk), .rst(phi_40_rst),
		.data_in_bus({{3'b0, phi_40_in1_data}, phi_40_in3_data, phi_40_in2_data}), .valid_in_bus({phi_40_in1_valid, phi_40_in3_valid, phi_40_in2_valid}), .ready_in_bus({phi_40_in1_ready, phi_40_in3_ready, phi_40_in2_ready}), 
		.data_out_bus({phi_40_out1_data}), .valid_out_bus({phi_40_out1_valid}), .ready_out_bus({phi_40_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_15
		(.clk(cst_15_clk), .rst(cst_15_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_15_in1_valid}), .ready_in_bus({cst_15_in1_ready}), 
		.data_out_bus({cst_15_out1_data}), .valid_out_bus({cst_15_out1_valid}), .ready_out_bus({cst_15_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_41
		(.clk(shl_41_clk), .rst(shl_41_rst),
		.data_in_bus({shl_41_in2_data, shl_41_in1_data}), .valid_in_bus({shl_41_in2_valid, shl_41_in1_valid}), .ready_in_bus({shl_41_in2_ready, shl_41_in1_ready}), 
		.data_out_bus({shl_41_out1_data}), .valid_out_bus({shl_41_out1_valid}), .ready_out_bus({shl_41_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_42
		(.clk(add_42_clk), .rst(add_42_rst),
		.data_in_bus({add_42_in2_data, add_42_in1_data}), .valid_in_bus({add_42_in2_valid, add_42_in1_valid}), .ready_in_bus({add_42_in2_ready, add_42_in1_ready}), 
		.data_out_bus({add_42_out1_data}), .valid_out_bus({add_42_out1_valid}), .ready_out_bus({add_42_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_load_op_load_45
		(.clk(load_45_clk), .rst(load_45_rst),
		.data_in_bus({load_45_in1_data}), .address_in_bus({load_45_in2_data}), .valid_in_bus({load_45_in2_valid, load_45_in1_valid}), .ready_in_bus({load_45_in2_ready, load_45_in1_ready}), 
		.data_out_bus({load_45_out1_data}), .address_out_bus({load_45_out2_data}), .valid_out_bus({load_45_out2_valid, load_45_out1_valid}), .ready_out_bus({load_45_out2_ready, load_45_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block9
		(.clk(brCst_block9_clk), .rst(brCst_block9_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block9_in1_valid}), .ready_in_bus({brCst_block9_in1_ready}), 
		.data_out_bus({brCst_block9_out1_data}), .valid_out_bus({brCst_block9_out1_valid}), .ready_out_bus({brCst_block9_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_16
		(.clk(cst_16_clk), .rst(cst_16_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_16_in1_valid}), .ready_in_bus({cst_16_in1_ready}), 
		.data_out_bus({cst_16_out1_data}), .valid_out_bus({cst_16_out1_valid}), .ready_out_bus({cst_16_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n13
		(.clk(phi_n13_clk), .rst(phi_n13_rst),
		.data_in_bus({phi_n13_in2_data, phi_n13_in1_data}), .valid_in_bus({phi_n13_in2_valid, phi_n13_in1_valid}), .ready_in_bus({phi_n13_in2_ready, phi_n13_in1_ready}), 
		.data_out_bus({phi_n13_out1_data}), .valid_out_bus({phi_n13_out1_valid}), .ready_out_bus({phi_n13_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_6
		(.clk(fork_6_clk), .rst(fork_6_rst),
		.data_in_bus({fork_6_in1_data}), .valid_in_bus({fork_6_in1_valid}), .ready_in_bus({fork_6_in1_ready}), 
		.data_out_bus({fork_6_out2_data, fork_6_out1_data}), .valid_out_bus({fork_6_out2_valid, fork_6_out1_valid}), .ready_out_bus({fork_6_out2_ready, fork_6_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_27
		(.clk(fork_27_clk), .rst(fork_27_rst),
		.data_in_bus({fork_27_in1_data}), .valid_in_bus({fork_27_in1_valid}), .ready_in_bus({fork_27_in1_ready}), 
		.data_out_bus({fork_27_out2_data, fork_27_out1_data}), .valid_out_bus({fork_27_out2_valid, fork_27_out1_valid}), .ready_out_bus({fork_27_out2_ready, fork_27_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_17
		(.clk(branch_17_clk), .rst(branch_17_rst),
		.data_in_bus({{31'b0, branch_17_in2_data}, branch_17_in1_data}), .valid_in_bus({branch_17_in2_valid, branch_17_in1_valid}), .ready_in_bus({branch_17_in2_ready, branch_17_in1_ready}), 
		.data_out_bus({branch_17_out2_data, branch_17_out1_data}), .valid_out_bus({branch_17_out2_valid, branch_17_out1_valid}), .ready_out_bus({branch_17_out2_ready, branch_17_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_18
		(.clk(branch_18_clk), .rst(branch_18_rst),
		.data_in_bus({{branch_18_in2_data}, branch_18_in1_data}), .valid_in_bus({branch_18_in2_valid, branch_18_in1_valid}), .ready_in_bus({branch_18_in2_ready, branch_18_in1_ready}), 
		.data_out_bus({branch_18_out2_data, branch_18_out1_data}), .valid_out_bus({branch_18_out2_valid, branch_18_out1_valid}), .ready_out_bus({branch_18_out2_ready, branch_18_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_19
		(.clk(branch_19_clk), .rst(branch_19_rst),
		.data_in_bus({{3'b0, branch_19_in2_data}, branch_19_in1_data}), .valid_in_bus({branch_19_in2_valid, branch_19_in1_valid}), .ready_in_bus({branch_19_in2_ready, branch_19_in1_ready}), 
		.data_out_bus({branch_19_out2_data, branch_19_out1_data}), .valid_out_bus({branch_19_out2_valid, branch_19_out1_valid}), .ready_out_bus({branch_19_out2_ready, branch_19_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_20
		(.clk(branch_20_clk), .rst(branch_20_rst),
		.data_in_bus({{3'b0, branch_20_in2_data}, branch_20_in1_data}), .valid_in_bus({branch_20_in2_valid, branch_20_in1_valid}), .ready_in_bus({branch_20_in2_ready, branch_20_in1_ready}), 
		.data_out_bus({branch_20_out2_data, branch_20_out1_data}), .valid_out_bus({branch_20_out2_valid, branch_20_out1_valid}), .ready_out_bus({branch_20_out2_ready, branch_20_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_41
		(.clk(fork_41_clk), .rst(fork_41_rst),
		.data_in_bus({fork_41_in1_data}), .valid_in_bus({fork_41_in1_valid}), .ready_in_bus({fork_41_in1_ready}), 
		.data_out_bus({fork_41_out5_data, fork_41_out4_data, fork_41_out3_data, fork_41_out2_data, fork_41_out1_data}), .valid_out_bus({fork_41_out5_valid, fork_41_out4_valid, fork_41_out3_valid, fork_41_out2_valid, fork_41_out1_valid}), .ready_out_bus({fork_41_out5_ready, fork_41_out4_ready, fork_41_out3_ready, fork_41_out2_ready, fork_41_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_28
		(.clk(phiC_28_clk), .rst(phiC_28_rst),
		.data_in_bus({phiC_28_in2_data, phiC_28_in1_data}), .valid_in_bus({phiC_28_in2_valid, phiC_28_in1_valid}), .ready_in_bus({phiC_28_in2_ready, phiC_28_in1_ready}), 
		.data_out_bus({phiC_28_out2_data, phiC_28_out1_data}), .valid_out_bus({phiC_28_out2_valid, phiC_28_out1_valid}), .ready_out_bus({phiC_28_out2_ready, phiC_28_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_63
		(.clk(forkC_63_clk), .rst(forkC_63_rst),
		.data_in_bus({forkC_63_in1_data}), .valid_in_bus({forkC_63_in1_valid}), .ready_in_bus({forkC_63_in1_ready}), 
		.data_out_bus({forkC_63_out3_data, forkC_63_out2_data, forkC_63_out1_data}), .valid_out_bus({forkC_63_out3_valid, forkC_63_out2_valid, forkC_63_out1_valid}), .ready_out_bus({forkC_63_out3_ready, forkC_63_out2_ready, forkC_63_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_50
		(.clk(branchC_50_clk), .rst(branchC_50_rst),
		.data_in_bus({{branchC_50_in2_data}, branchC_50_in1_data}), .valid_in_bus({branchC_50_in2_valid, branchC_50_in1_valid}), .ready_in_bus({branchC_50_in2_ready, branchC_50_in1_ready}), 
		.data_out_bus({branchC_50_out2_data, branchC_50_out1_data}), .valid_out_bus({branchC_50_out2_valid, branchC_50_out1_valid}), .ready_out_bus({branchC_50_out2_ready, branchC_50_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_10
		(.clk(source_10_clk), .rst(source_10_rst),
		.data_out_bus({source_10_out1_data}), .valid_out_bus({source_10_out1_valid}), .ready_out_bus({source_10_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block7
		(.clk(brCst_block7_clk), .rst(brCst_block7_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block7_in1_valid}), .ready_in_bus({brCst_block7_in1_ready}), 
		.data_out_bus({brCst_block7_out1_data}), .valid_out_bus({brCst_block7_out1_valid}), .ready_out_bus({brCst_block7_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_13
		(.clk(cst_13_clk), .rst(cst_13_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_13_in1_valid}), .ready_in_bus({cst_13_in1_ready}), 
		.data_out_bus({cst_13_out1_data}), .valid_out_bus({cst_13_out1_valid}), .ready_out_bus({cst_13_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_14
		(.clk(branch_14_clk), .rst(branch_14_rst),
		.data_in_bus({{branch_14_in2_data}, branch_14_in1_data}), .valid_in_bus({branch_14_in2_valid, branch_14_in1_valid}), .ready_in_bus({branch_14_in2_ready, branch_14_in1_ready}), 
		.data_out_bus({branch_14_out2_data, branch_14_out1_data}), .valid_out_bus({branch_14_out2_valid, branch_14_out1_valid}), .ready_out_bus({branch_14_out2_ready, branch_14_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_26
		(.clk(phiC_26_clk), .rst(phiC_26_rst),
		.data_in_bus({phiC_26_in1_data}), .valid_in_bus({phiC_26_in1_valid}), .ready_in_bus({phiC_26_in1_ready}), 
		.data_out_bus({phiC_26_out1_data}), .valid_out_bus({phiC_26_out1_valid}), .ready_out_bus({phiC_26_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_60
		(.clk(forkC_60_clk), .rst(forkC_60_rst),
		.data_in_bus({forkC_60_in1_data}), .valid_in_bus({forkC_60_in1_valid}), .ready_in_bus({forkC_60_in1_ready}), 
		.data_out_bus({forkC_60_out3_data, forkC_60_out2_data, forkC_60_out1_data}), .valid_out_bus({forkC_60_out3_valid, forkC_60_out2_valid, forkC_60_out1_valid}), .ready_out_bus({forkC_60_out3_ready, forkC_60_out2_ready, forkC_60_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_48
		(.clk(branchC_48_clk), .rst(branchC_48_rst),
		.data_in_bus({{branchC_48_in2_data}, branchC_48_in1_data}), .valid_in_bus({branchC_48_in2_valid, branchC_48_in1_valid}), .ready_in_bus({branchC_48_in2_ready, branchC_48_in1_ready}), 
		.data_out_bus({branchC_48_out2_data, branchC_48_out1_data}), .valid_out_bus({branchC_48_out2_valid, branchC_48_out1_valid}), .ready_out_bus({branchC_48_out2_ready, branchC_48_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_61
		(.clk(fork_61_clk), .rst(fork_61_rst),
		.data_in_bus({fork_61_in1_data}), .valid_in_bus({fork_61_in1_valid}), .ready_in_bus({fork_61_in1_ready}), 
		.data_out_bus({fork_61_out2_data, fork_61_out1_data}), .valid_out_bus({fork_61_out2_valid, fork_61_out1_valid}), .ready_out_bus({fork_61_out2_ready, fork_61_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block13
		(.clk(brCst_block13_clk), .rst(brCst_block13_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block13_in1_valid}), .ready_in_bus({brCst_block13_in1_ready}), 
		.data_out_bus({brCst_block13_out1_data}), .valid_out_bus({brCst_block13_out1_valid}), .ready_out_bus({brCst_block13_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_26
		(.clk(cst_26_clk), .rst(cst_26_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_26_in1_valid}), .ready_in_bus({cst_26_in1_ready}), 
		.data_out_bus({cst_26_out1_data}), .valid_out_bus({cst_26_out1_valid}), .ready_out_bus({cst_26_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_28
		(.clk(branch_28_clk), .rst(branch_28_rst),
		.data_in_bus({{branch_28_in2_data}, branch_28_in1_data}), .valid_in_bus({branch_28_in2_valid, branch_28_in1_valid}), .ready_in_bus({branch_28_in2_ready, branch_28_in1_ready}), 
		.data_out_bus({branch_28_out2_data, branch_28_out1_data}), .valid_out_bus({branch_28_out2_valid, branch_28_out1_valid}), .ready_out_bus({branch_28_out2_ready, branch_28_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_32
		(.clk(phiC_32_clk), .rst(phiC_32_rst),
		.data_in_bus({phiC_32_in1_data}), .valid_in_bus({phiC_32_in1_valid}), .ready_in_bus({phiC_32_in1_ready}), 
		.data_out_bus({phiC_32_out1_data}), .valid_out_bus({phiC_32_out1_valid}), .ready_out_bus({phiC_32_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_68
		(.clk(forkC_68_clk), .rst(forkC_68_rst),
		.data_in_bus({forkC_68_in1_data}), .valid_in_bus({forkC_68_in1_valid}), .ready_in_bus({forkC_68_in1_ready}), 
		.data_out_bus({forkC_68_out3_data, forkC_68_out2_data, forkC_68_out1_data}), .valid_out_bus({forkC_68_out3_valid, forkC_68_out2_valid, forkC_68_out1_valid}), .ready_out_bus({forkC_68_out3_ready, forkC_68_out2_ready, forkC_68_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_54
		(.clk(branchC_54_clk), .rst(branchC_54_rst),
		.data_in_bus({{branchC_54_in2_data}, branchC_54_in1_data}), .valid_in_bus({branchC_54_in2_valid, branchC_54_in1_valid}), .ready_in_bus({branchC_54_in2_ready, branchC_54_in1_ready}), 
		.data_out_bus({branchC_54_out2_data, branchC_54_out1_data}), .valid_out_bus({branchC_54_out2_valid, branchC_54_out1_valid}), .ready_out_bus({branchC_54_out2_ready, branchC_54_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_69
		(.clk(fork_69_clk), .rst(fork_69_rst),
		.data_in_bus({fork_69_in1_data}), .valid_in_bus({fork_69_in1_valid}), .ready_in_bus({fork_69_in1_ready}), 
		.data_out_bus({fork_69_out2_data, fork_69_out1_data}), .valid_out_bus({fork_69_out2_valid, fork_69_out1_valid}), .ready_out_bus({fork_69_out2_ready, fork_69_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4), .COND_SIZE(1)) mux_node_phi_75
		(.clk(phi_75_clk), .rst(phi_75_rst),
		.data_in_bus({{3'b0, phi_75_in1_data}, phi_75_in3_data, phi_75_in2_data}), .valid_in_bus({phi_75_in1_valid, phi_75_in3_valid, phi_75_in2_valid}), .ready_in_bus({phi_75_in1_ready, phi_75_in3_ready, phi_75_in2_ready}), 
		.data_out_bus({phi_75_out1_data}), .valid_out_bus({phi_75_out1_valid}), .ready_out_bus({phi_75_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block14
		(.clk(brCst_block14_clk), .rst(brCst_block14_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block14_in1_valid}), .ready_in_bus({brCst_block14_in1_ready}), 
		.data_out_bus({brCst_block14_out1_data}), .valid_out_bus({brCst_block14_out1_valid}), .ready_out_bus({brCst_block14_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_27
		(.clk(cst_27_clk), .rst(cst_27_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_27_in1_valid}), .ready_in_bus({cst_27_in1_ready}), 
		.data_out_bus({cst_27_out1_data}), .valid_out_bus({cst_27_out1_valid}), .ready_out_bus({cst_27_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_29
		(.clk(branch_29_clk), .rst(branch_29_rst),
		.data_in_bus({{branch_29_in2_data}, branch_29_in1_data}), .valid_in_bus({branch_29_in2_valid, branch_29_in1_valid}), .ready_in_bus({branch_29_in2_ready, branch_29_in1_ready}), 
		.data_out_bus({branch_29_out2_data, branch_29_out1_data}), .valid_out_bus({branch_29_out2_valid, branch_29_out1_valid}), .ready_out_bus({branch_29_out2_ready, branch_29_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_30
		(.clk(branch_30_clk), .rst(branch_30_rst),
		.data_in_bus({{3'b0, branch_30_in2_data}, branch_30_in1_data}), .valid_in_bus({branch_30_in2_valid, branch_30_in1_valid}), .ready_in_bus({branch_30_in2_ready, branch_30_in1_ready}), 
		.data_out_bus({branch_30_out2_data, branch_30_out1_data}), .valid_out_bus({branch_30_out2_valid, branch_30_out1_valid}), .ready_out_bus({branch_30_out2_ready, branch_30_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_46
		(.clk(fork_46_clk), .rst(fork_46_rst),
		.data_in_bus({fork_46_in1_data}), .valid_in_bus({fork_46_in1_valid}), .ready_in_bus({fork_46_in1_ready}), 
		.data_out_bus({fork_46_out3_data, fork_46_out2_data, fork_46_out1_data}), .valid_out_bus({fork_46_out3_valid, fork_46_out2_valid, fork_46_out1_valid}), .ready_out_bus({fork_46_out3_ready, fork_46_out2_ready, fork_46_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_33
		(.clk(phiC_33_clk), .rst(phiC_33_rst),
		.data_in_bus({phiC_33_in2_data, phiC_33_in1_data}), .valid_in_bus({phiC_33_in2_valid, phiC_33_in1_valid}), .ready_in_bus({phiC_33_in2_ready, phiC_33_in1_ready}), 
		.data_out_bus({phiC_33_out2_data, phiC_33_out1_data}), .valid_out_bus({phiC_33_out2_valid, phiC_33_out1_valid}), .ready_out_bus({phiC_33_out2_ready, phiC_33_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_70
		(.clk(forkC_70_clk), .rst(forkC_70_rst),
		.data_in_bus({forkC_70_in1_data}), .valid_in_bus({forkC_70_in1_valid}), .ready_in_bus({forkC_70_in1_ready}), 
		.data_out_bus({forkC_70_out3_data, forkC_70_out2_data, forkC_70_out1_data}), .valid_out_bus({forkC_70_out3_valid, forkC_70_out2_valid, forkC_70_out1_valid}), .ready_out_bus({forkC_70_out3_ready, forkC_70_out2_ready, forkC_70_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_55
		(.clk(branchC_55_clk), .rst(branchC_55_rst),
		.data_in_bus({{branchC_55_in2_data}, branchC_55_in1_data}), .valid_in_bus({branchC_55_in2_valid, branchC_55_in1_valid}), .ready_in_bus({branchC_55_in2_ready, branchC_55_in1_ready}), 
		.data_out_bus({branchC_55_out2_data, branchC_55_out1_data}), .valid_out_bus({branchC_55_out2_valid, branchC_55_out1_valid}), .ready_out_bus({branchC_55_out2_ready, branchC_55_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_37
		(.clk(cst_37_clk), .rst(cst_37_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_37_in1_valid}), .ready_in_bus({cst_37_in1_ready}), 
		.data_out_bus({cst_37_out1_data}), .valid_out_bus({cst_37_out1_valid}), .ready_out_bus({cst_37_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) add_op_add_108
		(.clk(add_108_clk), .rst(add_108_rst),
		.data_in_bus({add_108_in2_data, add_108_in1_data}), .valid_in_bus({add_108_in2_valid, add_108_in1_valid}), .ready_in_bus({add_108_in2_ready, add_108_in1_ready}), 
		.data_out_bus({add_108_out1_data}), .valid_out_bus({add_108_out1_valid}), .ready_out_bus({add_108_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) const_node_cst_38
		(.clk(cst_38_clk), .rst(cst_38_rst),
		.data_in_bus({4'd8}), .valid_in_bus({cst_38_in1_valid}), .ready_in_bus({cst_38_in1_ready}), 
		.data_out_bus({cst_38_out1_data}), .valid_out_bus({cst_38_out1_valid}), .ready_out_bus({cst_38_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_109
		(.clk(icmp_109_clk), .rst(icmp_109_rst),
		.data_in_bus({icmp_109_in2_data, icmp_109_in1_data}), .valid_in_bus({icmp_109_in2_valid, icmp_109_in1_valid}), .ready_in_bus({icmp_109_in2_ready, icmp_109_in1_ready}), 
		.data_out_bus({icmp_109_out1_data}), .valid_out_bus({icmp_109_out1_valid}), .ready_out_bus({icmp_109_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n14
		(.clk(phi_n14_clk), .rst(phi_n14_rst),
		.data_in_bus({phi_n14_in1_data}), .valid_in_bus({phi_n14_in1_valid}), .ready_in_bus({phi_n14_in1_ready}), 
		.data_out_bus({phi_n14_out1_data}), .valid_out_bus({phi_n14_out1_valid}), .ready_out_bus({phi_n14_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_17
		(.clk(fork_17_clk), .rst(fork_17_rst),
		.data_in_bus({fork_17_in1_data}), .valid_in_bus({fork_17_in1_valid}), .ready_in_bus({fork_17_in1_ready}), 
		.data_out_bus({fork_17_out2_data, fork_17_out1_data}), .valid_out_bus({fork_17_out2_valid, fork_17_out1_valid}), .ready_out_bus({fork_17_out2_ready, fork_17_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_41
		(.clk(branch_41_clk), .rst(branch_41_rst),
		.data_in_bus({{3'b0, branch_41_in2_data}, branch_41_in1_data}), .valid_in_bus({branch_41_in2_valid, branch_41_in1_valid}), .ready_in_bus({branch_41_in2_ready, branch_41_in1_ready}), 
		.data_out_bus({branch_41_out2_data, branch_41_out1_data}), .valid_out_bus({branch_41_out2_valid, branch_41_out1_valid}), .ready_out_bus({branch_41_out2_ready, branch_41_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_37
		(.clk(phiC_37_clk), .rst(phiC_37_rst),
		.data_in_bus({phiC_37_in1_data}), .valid_in_bus({phiC_37_in1_valid}), .ready_in_bus({phiC_37_in1_ready}), 
		.data_out_bus({phiC_37_out1_data}), .valid_out_bus({phiC_37_out1_valid}), .ready_out_bus({phiC_37_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_59
		(.clk(branchC_59_clk), .rst(branchC_59_rst),
		.data_in_bus({{branchC_59_in2_data}, branchC_59_in1_data}), .valid_in_bus({branchC_59_in2_valid, branchC_59_in1_valid}), .ready_in_bus({branchC_59_in2_ready, branchC_59_in1_ready}), 
		.data_out_bus({branchC_59_out2_data, branchC_59_out1_data}), .valid_out_bus({branchC_59_out2_valid, branchC_59_out1_valid}), .ready_out_bus({branchC_59_out2_ready, branchC_59_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_75
		(.clk(fork_75_clk), .rst(fork_75_rst),
		.data_in_bus({fork_75_in1_data}), .valid_in_bus({fork_75_in1_valid}), .ready_in_bus({fork_75_in1_ready}), 
		.data_out_bus({fork_75_out2_data, fork_75_out1_data}), .valid_out_bus({fork_75_out2_valid, fork_75_out1_valid}), .ready_out_bus({fork_75_out2_ready, fork_75_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_28
		(.clk(source_28_clk), .rst(source_28_rst),
		.data_out_bus({source_28_out1_data}), .valid_out_bus({source_28_out1_valid}), .ready_out_bus({source_28_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(4))source_node_source_29
		(.clk(source_29_clk), .rst(source_29_rst),
		.data_out_bus({source_29_out1_data}), .valid_out_bus({source_29_out1_valid}), .ready_out_bus({source_29_out1_ready}));

	ret_op #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) ret_op_ret_0
		(.clk(ret_0_clk), .rst(ret_0_rst),
		.data_in_bus({ret_0_in1_data}), .valid_in_bus({ret_0_in1_valid}), .ready_in_bus({ret_0_in1_ready}), 
		.data_out_bus({ret_0_out1_data}), .valid_out_bus({ret_0_out1_valid}), .ready_out_bus({ret_0_out1_ready}));

	end_node #(.INPUTS(1), .OUTPUTS(1), .MEMORY_INPUTS(7), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) end_node_end_0
		(.clk(end_0_clk), .rst(end_0_rst),
		.data_in_bus({end_0_in8_data}), .valid_in_bus({end_0_in8_valid}), .ready_in_bus({end_0_in8_ready}), .e_valid_bus({end_0_in7_valid, end_0_in6_valid, end_0_in5_valid, end_0_in4_valid, end_0_in3_valid, end_0_in2_valid, end_0_in1_valid}), .e_ready_bus({end_0_in7_ready, end_0_in6_ready, end_0_in5_ready, end_0_in4_ready, end_0_in3_ready, end_0_in2_ready, end_0_in1_ready}), 
		.data_out_bus({end_0_out1_data}), .valid_out_bus({end_0_out1_valid}), .ready_out_bus({end_0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_38
		(.clk(phiC_38_clk), .rst(phiC_38_rst),
		.data_in_bus({phiC_38_in1_data}), .valid_in_bus({phiC_38_in1_valid}), .ready_in_bus({phiC_38_in1_ready}), 
		.data_out_bus({phiC_38_out1_data}), .valid_out_bus({phiC_38_out1_valid}), .ready_out_bus({phiC_38_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_24
		(.clk(cst_24_clk), .rst(cst_24_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_24_in1_valid}), .ready_in_bus({cst_24_in1_ready}), 
		.data_out_bus({cst_24_out1_data}), .valid_out_bus({cst_24_out1_valid}), .ready_out_bus({cst_24_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) add_op_add_71
		(.clk(add_71_clk), .rst(add_71_rst),
		.data_in_bus({add_71_in2_data, add_71_in1_data}), .valid_in_bus({add_71_in2_valid, add_71_in1_valid}), .ready_in_bus({add_71_in2_ready, add_71_in1_ready}), 
		.data_out_bus({add_71_out1_data}), .valid_out_bus({add_71_out1_valid}), .ready_out_bus({add_71_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) const_node_cst_25
		(.clk(cst_25_clk), .rst(cst_25_rst),
		.data_in_bus({4'd8}), .valid_in_bus({cst_25_in1_valid}), .ready_in_bus({cst_25_in1_ready}), 
		.data_out_bus({cst_25_out1_data}), .valid_out_bus({cst_25_out1_valid}), .ready_out_bus({cst_25_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_72
		(.clk(icmp_72_clk), .rst(icmp_72_rst),
		.data_in_bus({icmp_72_in2_data, icmp_72_in1_data}), .valid_in_bus({icmp_72_in2_valid, icmp_72_in1_valid}), .ready_in_bus({icmp_72_in2_ready, icmp_72_in1_ready}), 
		.data_out_bus({icmp_72_out1_data}), .valid_out_bus({icmp_72_out1_valid}), .ready_out_bus({icmp_72_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n12
		(.clk(phi_n12_clk), .rst(phi_n12_rst),
		.data_in_bus({phi_n12_in1_data}), .valid_in_bus({phi_n12_in1_valid}), .ready_in_bus({phi_n12_in1_ready}), 
		.data_out_bus({phi_n12_out1_data}), .valid_out_bus({phi_n12_out1_valid}), .ready_out_bus({phi_n12_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_11
		(.clk(fork_11_clk), .rst(fork_11_rst),
		.data_in_bus({fork_11_in1_data}), .valid_in_bus({fork_11_in1_valid}), .ready_in_bus({fork_11_in1_ready}), 
		.data_out_bus({fork_11_out2_data, fork_11_out1_data}), .valid_out_bus({fork_11_out2_valid, fork_11_out1_valid}), .ready_out_bus({fork_11_out2_ready, fork_11_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_27
		(.clk(branch_27_clk), .rst(branch_27_rst),
		.data_in_bus({{3'b0, branch_27_in2_data}, branch_27_in1_data}), .valid_in_bus({branch_27_in2_valid, branch_27_in1_valid}), .ready_in_bus({branch_27_in2_ready, branch_27_in1_ready}), 
		.data_out_bus({branch_27_out2_data, branch_27_out1_data}), .valid_out_bus({branch_27_out2_valid, branch_27_out1_valid}), .ready_out_bus({branch_27_out2_ready, branch_27_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_31
		(.clk(phiC_31_clk), .rst(phiC_31_rst),
		.data_in_bus({phiC_31_in1_data}), .valid_in_bus({phiC_31_in1_valid}), .ready_in_bus({phiC_31_in1_ready}), 
		.data_out_bus({phiC_31_out1_data}), .valid_out_bus({phiC_31_out1_valid}), .ready_out_bus({phiC_31_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_53
		(.clk(branchC_53_clk), .rst(branchC_53_rst),
		.data_in_bus({{branchC_53_in2_data}, branchC_53_in1_data}), .valid_in_bus({branchC_53_in2_valid, branchC_53_in1_valid}), .ready_in_bus({branchC_53_in2_ready, branchC_53_in1_ready}), 
		.data_out_bus({branchC_53_out2_data, branchC_53_out1_data}), .valid_out_bus({branchC_53_out2_valid, branchC_53_out1_valid}), .ready_out_bus({branchC_53_out2_ready, branchC_53_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_67
		(.clk(fork_67_clk), .rst(fork_67_rst),
		.data_in_bus({fork_67_in1_data}), .valid_in_bus({fork_67_in1_valid}), .ready_in_bus({fork_67_in1_ready}), 
		.data_out_bus({fork_67_out2_data, fork_67_out1_data}), .valid_out_bus({fork_67_out2_valid, fork_67_out1_valid}), .ready_out_bus({fork_67_out2_ready, fork_67_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_18
		(.clk(source_18_clk), .rst(source_18_rst),
		.data_out_bus({source_18_out1_data}), .valid_out_bus({source_18_out1_valid}), .ready_out_bus({source_18_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(4))source_node_source_19
		(.clk(source_19_clk), .rst(source_19_rst),
		.data_out_bus({source_19_out1_data}), .valid_out_bus({source_19_out1_valid}), .ready_out_bus({source_19_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_47
		(.clk(phi_47_clk), .rst(phi_47_rst),
		.data_in_bus({{31'b0, phi_47_in1_data}, phi_47_in3_data, phi_47_in2_data}), .valid_in_bus({phi_47_in1_valid, phi_47_in3_valid, phi_47_in2_valid}), .ready_in_bus({phi_47_in1_ready, phi_47_in3_ready, phi_47_in2_ready}), 
		.data_out_bus({phi_47_out1_data}), .valid_out_bus({phi_47_out1_valid}), .ready_out_bus({phi_47_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4), .COND_SIZE(1)) mux_node_phi_48
		(.clk(phi_48_clk), .rst(phi_48_rst),
		.data_in_bus({{3'b0, phi_48_in1_data}, phi_48_in3_data, phi_48_in2_data}), .valid_in_bus({phi_48_in1_valid, phi_48_in3_valid, phi_48_in2_valid}), .ready_in_bus({phi_48_in1_ready, phi_48_in3_ready, phi_48_in2_ready}), 
		.data_out_bus({phi_48_out1_data}), .valid_out_bus({phi_48_out1_valid}), .ready_out_bus({phi_48_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_17
		(.clk(cst_17_clk), .rst(cst_17_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_17_in1_valid}), .ready_in_bus({cst_17_in1_ready}), 
		.data_out_bus({cst_17_out1_data}), .valid_out_bus({cst_17_out1_valid}), .ready_out_bus({cst_17_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_49
		(.clk(shl_49_clk), .rst(shl_49_rst),
		.data_in_bus({shl_49_in2_data, shl_49_in1_data}), .valid_in_bus({shl_49_in2_valid, shl_49_in1_valid}), .ready_in_bus({shl_49_in2_ready, shl_49_in1_ready}), 
		.data_out_bus({shl_49_out1_data}), .valid_out_bus({shl_49_out1_valid}), .ready_out_bus({shl_49_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_50
		(.clk(add_50_clk), .rst(add_50_rst),
		.data_in_bus({add_50_in2_data, add_50_in1_data}), .valid_in_bus({add_50_in2_valid, add_50_in1_valid}), .ready_in_bus({add_50_in2_ready, add_50_in1_ready}), 
		.data_out_bus({add_50_out1_data}), .valid_out_bus({add_50_out1_valid}), .ready_out_bus({add_50_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_load_op_load_53
		(.clk(load_53_clk), .rst(load_53_rst),
		.data_in_bus({load_53_in1_data}), .address_in_bus({load_53_in2_data}), .valid_in_bus({load_53_in2_valid, load_53_in1_valid}), .ready_in_bus({load_53_in2_ready, load_53_in1_ready}), 
		.data_out_bus({load_53_out1_data}), .address_out_bus({load_53_out2_data}), .valid_out_bus({load_53_out2_valid, load_53_out1_valid}), .ready_out_bus({load_53_out2_ready, load_53_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_18
		(.clk(cst_18_clk), .rst(cst_18_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_18_in1_valid}), .ready_in_bus({cst_18_in1_ready}), 
		.data_out_bus({cst_18_out1_data}), .valid_out_bus({cst_18_out1_valid}), .ready_out_bus({cst_18_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_54
		(.clk(shl_54_clk), .rst(shl_54_rst),
		.data_in_bus({shl_54_in2_data, shl_54_in1_data}), .valid_in_bus({shl_54_in2_valid, shl_54_in1_valid}), .ready_in_bus({shl_54_in2_ready, shl_54_in1_ready}), 
		.data_out_bus({shl_54_out1_data}), .valid_out_bus({shl_54_out1_valid}), .ready_out_bus({shl_54_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_55
		(.clk(add_55_clk), .rst(add_55_rst),
		.data_in_bus({add_55_in2_data, add_55_in1_data}), .valid_in_bus({add_55_in2_valid, add_55_in1_valid}), .ready_in_bus({add_55_in2_ready, add_55_in1_ready}), 
		.data_out_bus({add_55_out1_data}), .valid_out_bus({add_55_out1_valid}), .ready_out_bus({add_55_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_load_op_load_58
		(.clk(load_58_clk), .rst(load_58_rst),
		.data_in_bus({load_58_in1_data}), .address_in_bus({load_58_in2_data}), .valid_in_bus({load_58_in2_valid, load_58_in1_valid}), .ready_in_bus({load_58_in2_ready, load_58_in1_ready}), 
		.data_out_bus({load_58_out1_data}), .address_out_bus({load_58_out2_data}), .valid_out_bus({load_58_out2_valid, load_58_out1_valid}), .ready_out_bus({load_58_out2_ready, load_58_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_19
		(.clk(cst_19_clk), .rst(cst_19_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_19_in1_valid}), .ready_in_bus({cst_19_in1_ready}), 
		.data_out_bus({cst_19_out1_data}), .valid_out_bus({cst_19_out1_valid}), .ready_out_bus({cst_19_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) add_op_add_61
		(.clk(add_61_clk), .rst(add_61_rst),
		.data_in_bus({add_61_in2_data, add_61_in1_data}), .valid_in_bus({add_61_in2_valid, add_61_in1_valid}), .ready_in_bus({add_61_in2_ready, add_61_in1_ready}), 
		.data_out_bus({add_61_out1_data}), .valid_out_bus({add_61_out1_valid}), .ready_out_bus({add_61_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) const_node_cst_20
		(.clk(cst_20_clk), .rst(cst_20_rst),
		.data_in_bus({4'd8}), .valid_in_bus({cst_20_in1_valid}), .ready_in_bus({cst_20_in1_ready}), 
		.data_out_bus({cst_20_out1_data}), .valid_out_bus({cst_20_out1_valid}), .ready_out_bus({cst_20_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_62
		(.clk(icmp_62_clk), .rst(icmp_62_rst),
		.data_in_bus({icmp_62_in2_data, icmp_62_in1_data}), .valid_in_bus({icmp_62_in2_valid, icmp_62_in1_valid}), .ready_in_bus({icmp_62_in2_ready, icmp_62_in1_ready}), 
		.data_out_bus({icmp_62_out1_data}), .valid_out_bus({icmp_62_out1_valid}), .ready_out_bus({icmp_62_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n10
		(.clk(phi_n10_clk), .rst(phi_n10_rst),
		.data_in_bus({phi_n10_in2_data, phi_n10_in1_data}), .valid_in_bus({phi_n10_in2_valid, phi_n10_in1_valid}), .ready_in_bus({phi_n10_in2_ready, phi_n10_in1_ready}), 
		.data_out_bus({phi_n10_out1_data}), .valid_out_bus({phi_n10_out1_valid}), .ready_out_bus({phi_n10_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n11
		(.clk(phi_n11_clk), .rst(phi_n11_rst),
		.data_in_bus({phi_n11_in2_data, phi_n11_in1_data}), .valid_in_bus({phi_n11_in2_valid, phi_n11_in1_valid}), .ready_in_bus({phi_n11_in2_ready, phi_n11_in1_ready}), 
		.data_out_bus({phi_n11_out1_data}), .valid_out_bus({phi_n11_out1_valid}), .ready_out_bus({phi_n11_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_7
		(.clk(fork_7_clk), .rst(fork_7_rst),
		.data_in_bus({fork_7_in1_data}), .valid_in_bus({fork_7_in1_valid}), .ready_in_bus({fork_7_in1_ready}), 
		.data_out_bus({fork_7_out3_data, fork_7_out2_data, fork_7_out1_data}), .valid_out_bus({fork_7_out3_valid, fork_7_out2_valid, fork_7_out1_valid}), .ready_out_bus({fork_7_out3_ready, fork_7_out2_ready, fork_7_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_9
		(.clk(fork_9_clk), .rst(fork_9_rst),
		.data_in_bus({fork_9_in1_data}), .valid_in_bus({fork_9_in1_valid}), .ready_in_bus({fork_9_in1_ready}), 
		.data_out_bus({fork_9_out2_data, fork_9_out1_data}), .valid_out_bus({fork_9_out2_valid, fork_9_out1_valid}), .ready_out_bus({fork_9_out2_ready, fork_9_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_25
		(.clk(fork_25_clk), .rst(fork_25_rst),
		.data_in_bus({fork_25_in1_data}), .valid_in_bus({fork_25_in1_valid}), .ready_in_bus({fork_25_in1_ready}), 
		.data_out_bus({fork_25_out2_data, fork_25_out1_data}), .valid_out_bus({fork_25_out2_valid, fork_25_out1_valid}), .ready_out_bus({fork_25_out2_ready, fork_25_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_26
		(.clk(fork_26_clk), .rst(fork_26_rst),
		.data_in_bus({fork_26_in1_data}), .valid_in_bus({fork_26_in1_valid}), .ready_in_bus({fork_26_in1_ready}), 
		.data_out_bus({fork_26_out2_data, fork_26_out1_data}), .valid_out_bus({fork_26_out2_valid, fork_26_out1_valid}), .ready_out_bus({fork_26_out2_ready, fork_26_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_21
		(.clk(branch_21_clk), .rst(branch_21_rst),
		.data_in_bus({{31'b0, branch_21_in2_data}, branch_21_in1_data}), .valid_in_bus({branch_21_in2_valid, branch_21_in1_valid}), .ready_in_bus({branch_21_in2_ready, branch_21_in1_ready}), 
		.data_out_bus({branch_21_out2_data, branch_21_out1_data}), .valid_out_bus({branch_21_out2_valid, branch_21_out1_valid}), .ready_out_bus({branch_21_out2_ready, branch_21_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_22
		(.clk(branch_22_clk), .rst(branch_22_rst),
		.data_in_bus({{3'b0, branch_22_in2_data}, branch_22_in1_data}), .valid_in_bus({branch_22_in2_valid, branch_22_in1_valid}), .ready_in_bus({branch_22_in2_ready, branch_22_in1_ready}), 
		.data_out_bus({branch_22_out2_data, branch_22_out1_data}), .valid_out_bus({branch_22_out2_valid, branch_22_out1_valid}), .ready_out_bus({branch_22_out2_ready, branch_22_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_23
		(.clk(branch_23_clk), .rst(branch_23_rst),
		.data_in_bus({{3'b0, branch_23_in2_data}, branch_23_in1_data}), .valid_in_bus({branch_23_in2_valid, branch_23_in1_valid}), .ready_in_bus({branch_23_in2_ready, branch_23_in1_ready}), 
		.data_out_bus({branch_23_out2_data, branch_23_out1_data}), .valid_out_bus({branch_23_out2_valid, branch_23_out1_valid}), .ready_out_bus({branch_23_out2_ready, branch_23_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_24
		(.clk(branch_24_clk), .rst(branch_24_rst),
		.data_in_bus({{3'b0, branch_24_in2_data}, branch_24_in1_data}), .valid_in_bus({branch_24_in2_valid, branch_24_in1_valid}), .ready_in_bus({branch_24_in2_ready, branch_24_in1_ready}), 
		.data_out_bus({branch_24_out2_data, branch_24_out1_data}), .valid_out_bus({branch_24_out2_valid, branch_24_out1_valid}), .ready_out_bus({branch_24_out2_ready, branch_24_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_42
		(.clk(fork_42_clk), .rst(fork_42_rst),
		.data_in_bus({fork_42_in1_data}), .valid_in_bus({fork_42_in1_valid}), .ready_in_bus({fork_42_in1_ready}), 
		.data_out_bus({fork_42_out5_data, fork_42_out4_data, fork_42_out3_data, fork_42_out2_data, fork_42_out1_data}), .valid_out_bus({fork_42_out5_valid, fork_42_out4_valid, fork_42_out3_valid, fork_42_out2_valid, fork_42_out1_valid}), .ready_out_bus({fork_42_out5_ready, fork_42_out4_ready, fork_42_out3_ready, fork_42_out2_ready, fork_42_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_29
		(.clk(phiC_29_clk), .rst(phiC_29_rst),
		.data_in_bus({phiC_29_in2_data, phiC_29_in1_data}), .valid_in_bus({phiC_29_in2_valid, phiC_29_in1_valid}), .ready_in_bus({phiC_29_in2_ready, phiC_29_in1_ready}), 
		.data_out_bus({phiC_29_out2_data, phiC_29_out1_data}), .valid_out_bus({phiC_29_out2_valid, phiC_29_out1_valid}), .ready_out_bus({phiC_29_out2_ready, phiC_29_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_51
		(.clk(branchC_51_clk), .rst(branchC_51_rst),
		.data_in_bus({{branchC_51_in2_data}, branchC_51_in1_data}), .valid_in_bus({branchC_51_in2_valid, branchC_51_in1_valid}), .ready_in_bus({branchC_51_in2_ready, branchC_51_in1_ready}), 
		.data_out_bus({branchC_51_out2_data, branchC_51_out1_data}), .valid_out_bus({branchC_51_out2_valid, branchC_51_out1_valid}), .ready_out_bus({branchC_51_out2_ready, branchC_51_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_11
		(.clk(source_11_clk), .rst(source_11_rst),
		.data_out_bus({source_11_out1_data}), .valid_out_bus({source_11_out1_valid}), .ready_out_bus({source_11_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_12
		(.clk(source_12_clk), .rst(source_12_rst),
		.data_out_bus({source_12_out1_data}), .valid_out_bus({source_12_out1_valid}), .ready_out_bus({source_12_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_13
		(.clk(source_13_clk), .rst(source_13_rst),
		.data_out_bus({source_13_out1_data}), .valid_out_bus({source_13_out1_valid}), .ready_out_bus({source_13_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(4))source_node_source_14
		(.clk(source_14_clk), .rst(source_14_rst),
		.data_out_bus({source_14_out1_data}), .valid_out_bus({source_14_out1_valid}), .ready_out_bus({source_14_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_82
		(.clk(fork_82_clk), .rst(fork_82_rst),
		.data_in_bus({fork_82_in1_data}), .valid_in_bus({fork_82_in1_valid}), .ready_in_bus({fork_82_in1_ready}), 
		.data_out_bus({fork_82_out2_data, fork_82_out1_data}), .valid_out_bus({fork_82_out2_valid, fork_82_out1_valid}), .ready_out_bus({fork_82_out2_ready, fork_82_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_10
		(.clk(phi_10_clk), .rst(phi_10_rst),
		.data_in_bus({{31'b0, phi_10_in1_data}, phi_10_in3_data, phi_10_in2_data}), .valid_in_bus({phi_10_in1_valid, phi_10_in3_valid, phi_10_in2_valid}), .ready_in_bus({phi_10_in1_ready, phi_10_in3_ready, phi_10_in2_ready}), 
		.data_out_bus({phi_10_out1_data}), .valid_out_bus({phi_10_out1_valid}), .ready_out_bus({phi_10_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4), .COND_SIZE(1)) mux_node_phi_11
		(.clk(phi_11_clk), .rst(phi_11_rst),
		.data_in_bus({{3'b0, phi_11_in1_data}, phi_11_in3_data, phi_11_in2_data}), .valid_in_bus({phi_11_in1_valid, phi_11_in3_valid, phi_11_in2_valid}), .ready_in_bus({phi_11_in1_ready, phi_11_in3_ready, phi_11_in2_ready}), 
		.data_out_bus({phi_11_out1_data}), .valid_out_bus({phi_11_out1_valid}), .ready_out_bus({phi_11_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_4
		(.clk(cst_4_clk), .rst(cst_4_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_4_in1_valid}), .ready_in_bus({cst_4_in1_ready}), 
		.data_out_bus({cst_4_out1_data}), .valid_out_bus({cst_4_out1_valid}), .ready_out_bus({cst_4_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_12
		(.clk(shl_12_clk), .rst(shl_12_rst),
		.data_in_bus({shl_12_in2_data, shl_12_in1_data}), .valid_in_bus({shl_12_in2_valid, shl_12_in1_valid}), .ready_in_bus({shl_12_in2_ready, shl_12_in1_ready}), 
		.data_out_bus({shl_12_out1_data}), .valid_out_bus({shl_12_out1_valid}), .ready_out_bus({shl_12_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_13
		(.clk(add_13_clk), .rst(add_13_rst),
		.data_in_bus({add_13_in2_data, add_13_in1_data}), .valid_in_bus({add_13_in2_valid, add_13_in1_valid}), .ready_in_bus({add_13_in2_ready, add_13_in1_ready}), 
		.data_out_bus({add_13_out1_data}), .valid_out_bus({add_13_out1_valid}), .ready_out_bus({add_13_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_load_op_load_16
		(.clk(load_16_clk), .rst(load_16_rst),
		.data_in_bus({load_16_in1_data}), .address_in_bus({load_16_in2_data}), .valid_in_bus({load_16_in2_valid, load_16_in1_valid}), .ready_in_bus({load_16_in2_ready, load_16_in1_ready}), 
		.data_out_bus({load_16_out1_data}), .address_out_bus({load_16_out2_data}), .valid_out_bus({load_16_out2_valid, load_16_out1_valid}), .ready_out_bus({load_16_out2_ready, load_16_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_5
		(.clk(cst_5_clk), .rst(cst_5_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_5_in1_valid}), .ready_in_bus({cst_5_in1_ready}), 
		.data_out_bus({cst_5_out1_data}), .valid_out_bus({cst_5_out1_valid}), .ready_out_bus({cst_5_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_17
		(.clk(shl_17_clk), .rst(shl_17_rst),
		.data_in_bus({shl_17_in2_data, shl_17_in1_data}), .valid_in_bus({shl_17_in2_valid, shl_17_in1_valid}), .ready_in_bus({shl_17_in2_ready, shl_17_in1_ready}), 
		.data_out_bus({shl_17_out1_data}), .valid_out_bus({shl_17_out1_valid}), .ready_out_bus({shl_17_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_18
		(.clk(add_18_clk), .rst(add_18_rst),
		.data_in_bus({add_18_in2_data, add_18_in1_data}), .valid_in_bus({add_18_in2_valid, add_18_in1_valid}), .ready_in_bus({add_18_in2_ready, add_18_in1_ready}), 
		.data_out_bus({add_18_out1_data}), .valid_out_bus({add_18_out1_valid}), .ready_out_bus({add_18_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_load_op_load_21
		(.clk(load_21_clk), .rst(load_21_rst),
		.data_in_bus({load_21_in1_data}), .address_in_bus({load_21_in2_data}), .valid_in_bus({load_21_in2_valid, load_21_in1_valid}), .ready_in_bus({load_21_in2_ready, load_21_in1_ready}), 
		.data_out_bus({load_21_out1_data}), .address_out_bus({load_21_out2_data}), .valid_out_bus({load_21_out2_valid, load_21_out1_valid}), .ready_out_bus({load_21_out2_ready, load_21_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_6
		(.clk(cst_6_clk), .rst(cst_6_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_6_in1_valid}), .ready_in_bus({cst_6_in1_ready}), 
		.data_out_bus({cst_6_out1_data}), .valid_out_bus({cst_6_out1_valid}), .ready_out_bus({cst_6_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) add_op_add_24
		(.clk(add_24_clk), .rst(add_24_rst),
		.data_in_bus({add_24_in2_data, add_24_in1_data}), .valid_in_bus({add_24_in2_valid, add_24_in1_valid}), .ready_in_bus({add_24_in2_ready, add_24_in1_ready}), 
		.data_out_bus({add_24_out1_data}), .valid_out_bus({add_24_out1_valid}), .ready_out_bus({add_24_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) const_node_cst_7
		(.clk(cst_7_clk), .rst(cst_7_rst),
		.data_in_bus({4'd8}), .valid_in_bus({cst_7_in1_valid}), .ready_in_bus({cst_7_in1_ready}), 
		.data_out_bus({cst_7_out1_data}), .valid_out_bus({cst_7_out1_valid}), .ready_out_bus({cst_7_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_25
		(.clk(icmp_25_clk), .rst(icmp_25_rst),
		.data_in_bus({icmp_25_in2_data, icmp_25_in1_data}), .valid_in_bus({icmp_25_in2_valid, icmp_25_in1_valid}), .ready_in_bus({icmp_25_in2_ready, icmp_25_in1_ready}), 
		.data_out_bus({icmp_25_out1_data}), .valid_out_bus({icmp_25_out1_valid}), .ready_out_bus({icmp_25_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n8
		(.clk(phi_n8_clk), .rst(phi_n8_rst),
		.data_in_bus({phi_n8_in2_data, phi_n8_in1_data}), .valid_in_bus({phi_n8_in2_valid, phi_n8_in1_valid}), .ready_in_bus({phi_n8_in2_ready, phi_n8_in1_ready}), 
		.data_out_bus({phi_n8_out1_data}), .valid_out_bus({phi_n8_out1_valid}), .ready_out_bus({phi_n8_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n9
		(.clk(phi_n9_clk), .rst(phi_n9_rst),
		.data_in_bus({phi_n9_in2_data, phi_n9_in1_data}), .valid_in_bus({phi_n9_in2_valid, phi_n9_in1_valid}), .ready_in_bus({phi_n9_in2_ready, phi_n9_in1_ready}), 
		.data_out_bus({phi_n9_out1_data}), .valid_out_bus({phi_n9_out1_valid}), .ready_out_bus({phi_n9_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_1
		(.clk(fork_1_clk), .rst(fork_1_rst),
		.data_in_bus({fork_1_in1_data}), .valid_in_bus({fork_1_in1_valid}), .ready_in_bus({fork_1_in1_ready}), 
		.data_out_bus({fork_1_out3_data, fork_1_out2_data, fork_1_out1_data}), .valid_out_bus({fork_1_out3_valid, fork_1_out2_valid, fork_1_out1_valid}), .ready_out_bus({fork_1_out3_ready, fork_1_out2_ready, fork_1_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_3
		(.clk(fork_3_clk), .rst(fork_3_rst),
		.data_in_bus({fork_3_in1_data}), .valid_in_bus({fork_3_in1_valid}), .ready_in_bus({fork_3_in1_ready}), 
		.data_out_bus({fork_3_out2_data, fork_3_out1_data}), .valid_out_bus({fork_3_out2_valid, fork_3_out1_valid}), .ready_out_bus({fork_3_out2_ready, fork_3_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_23
		(.clk(fork_23_clk), .rst(fork_23_rst),
		.data_in_bus({fork_23_in1_data}), .valid_in_bus({fork_23_in1_valid}), .ready_in_bus({fork_23_in1_ready}), 
		.data_out_bus({fork_23_out2_data, fork_23_out1_data}), .valid_out_bus({fork_23_out2_valid, fork_23_out1_valid}), .ready_out_bus({fork_23_out2_ready, fork_23_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_24
		(.clk(fork_24_clk), .rst(fork_24_rst),
		.data_in_bus({fork_24_in1_data}), .valid_in_bus({fork_24_in1_valid}), .ready_in_bus({fork_24_in1_ready}), 
		.data_out_bus({fork_24_out2_data, fork_24_out1_data}), .valid_out_bus({fork_24_out2_valid, fork_24_out1_valid}), .ready_out_bus({fork_24_out2_ready, fork_24_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_7
		(.clk(branch_7_clk), .rst(branch_7_rst),
		.data_in_bus({{31'b0, branch_7_in2_data}, branch_7_in1_data}), .valid_in_bus({branch_7_in2_valid, branch_7_in1_valid}), .ready_in_bus({branch_7_in2_ready, branch_7_in1_ready}), 
		.data_out_bus({branch_7_out2_data, branch_7_out1_data}), .valid_out_bus({branch_7_out2_valid, branch_7_out1_valid}), .ready_out_bus({branch_7_out2_ready, branch_7_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_8
		(.clk(branch_8_clk), .rst(branch_8_rst),
		.data_in_bus({{3'b0, branch_8_in2_data}, branch_8_in1_data}), .valid_in_bus({branch_8_in2_valid, branch_8_in1_valid}), .ready_in_bus({branch_8_in2_ready, branch_8_in1_ready}), 
		.data_out_bus({branch_8_out2_data, branch_8_out1_data}), .valid_out_bus({branch_8_out2_valid, branch_8_out1_valid}), .ready_out_bus({branch_8_out2_ready, branch_8_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_9
		(.clk(branch_9_clk), .rst(branch_9_rst),
		.data_in_bus({{3'b0, branch_9_in2_data}, branch_9_in1_data}), .valid_in_bus({branch_9_in2_valid, branch_9_in1_valid}), .ready_in_bus({branch_9_in2_ready, branch_9_in1_ready}), 
		.data_out_bus({branch_9_out2_data, branch_9_out1_data}), .valid_out_bus({branch_9_out2_valid, branch_9_out1_valid}), .ready_out_bus({branch_9_out2_ready, branch_9_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_10
		(.clk(branch_10_clk), .rst(branch_10_rst),
		.data_in_bus({{3'b0, branch_10_in2_data}, branch_10_in1_data}), .valid_in_bus({branch_10_in2_valid, branch_10_in1_valid}), .ready_in_bus({branch_10_in2_ready, branch_10_in1_ready}), 
		.data_out_bus({branch_10_out2_data, branch_10_out1_data}), .valid_out_bus({branch_10_out2_valid, branch_10_out1_valid}), .ready_out_bus({branch_10_out2_ready, branch_10_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_36
		(.clk(fork_36_clk), .rst(fork_36_rst),
		.data_in_bus({fork_36_in1_data}), .valid_in_bus({fork_36_in1_valid}), .ready_in_bus({fork_36_in1_ready}), 
		.data_out_bus({fork_36_out5_data, fork_36_out4_data, fork_36_out3_data, fork_36_out2_data, fork_36_out1_data}), .valid_out_bus({fork_36_out5_valid, fork_36_out4_valid, fork_36_out3_valid, fork_36_out2_valid, fork_36_out1_valid}), .ready_out_bus({fork_36_out5_ready, fork_36_out4_ready, fork_36_out3_ready, fork_36_out2_ready, fork_36_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_23
		(.clk(phiC_23_clk), .rst(phiC_23_rst),
		.data_in_bus({phiC_23_in2_data, phiC_23_in1_data}), .valid_in_bus({phiC_23_in2_valid, phiC_23_in1_valid}), .ready_in_bus({phiC_23_in2_ready, phiC_23_in1_ready}), 
		.data_out_bus({phiC_23_out2_data, phiC_23_out1_data}), .valid_out_bus({phiC_23_out2_valid, phiC_23_out1_valid}), .ready_out_bus({phiC_23_out2_ready, phiC_23_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_45
		(.clk(branchC_45_clk), .rst(branchC_45_rst),
		.data_in_bus({{branchC_45_in2_data}, branchC_45_in1_data}), .valid_in_bus({branchC_45_in2_valid, branchC_45_in1_valid}), .ready_in_bus({branchC_45_in2_ready, branchC_45_in1_ready}), 
		.data_out_bus({branchC_45_out2_data, branchC_45_out1_data}), .valid_out_bus({branchC_45_out2_valid, branchC_45_out1_valid}), .ready_out_bus({branchC_45_out2_ready, branchC_45_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_1
		(.clk(source_1_clk), .rst(source_1_rst),
		.data_out_bus({source_1_out1_data}), .valid_out_bus({source_1_out1_valid}), .ready_out_bus({source_1_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_2
		(.clk(source_2_clk), .rst(source_2_rst),
		.data_out_bus({source_2_out1_data}), .valid_out_bus({source_2_out1_valid}), .ready_out_bus({source_2_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_3
		(.clk(source_3_clk), .rst(source_3_rst),
		.data_out_bus({source_3_out1_data}), .valid_out_bus({source_3_out1_valid}), .ready_out_bus({source_3_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(4))source_node_source_4
		(.clk(source_4_clk), .rst(source_4_rst),
		.data_out_bus({source_4_out1_data}), .valid_out_bus({source_4_out1_valid}), .ready_out_bus({source_4_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_79
		(.clk(fork_79_clk), .rst(fork_79_rst),
		.data_in_bus({fork_79_in1_data}), .valid_in_bus({fork_79_in1_valid}), .ready_in_bus({fork_79_in1_ready}), 
		.data_out_bus({fork_79_out2_data, fork_79_out1_data}), .valid_out_bus({fork_79_out2_valid, fork_79_out1_valid}), .ready_out_bus({fork_79_out2_ready, fork_79_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_84
		(.clk(phi_84_clk), .rst(phi_84_rst),
		.data_in_bus({{31'b0, phi_84_in1_data}, phi_84_in3_data, phi_84_in2_data}), .valid_in_bus({phi_84_in1_valid, phi_84_in3_valid, phi_84_in2_valid}), .ready_in_bus({phi_84_in1_ready, phi_84_in3_ready, phi_84_in2_ready}), 
		.data_out_bus({phi_84_out1_data}), .valid_out_bus({phi_84_out1_valid}), .ready_out_bus({phi_84_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4), .COND_SIZE(1)) mux_node_phi_85
		(.clk(phi_85_clk), .rst(phi_85_rst),
		.data_in_bus({{3'b0, phi_85_in1_data}, phi_85_in3_data, phi_85_in2_data}), .valid_in_bus({phi_85_in1_valid, phi_85_in3_valid, phi_85_in2_valid}), .ready_in_bus({phi_85_in1_ready, phi_85_in3_ready, phi_85_in2_ready}), 
		.data_out_bus({phi_85_out1_data}), .valid_out_bus({phi_85_out1_valid}), .ready_out_bus({phi_85_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_30
		(.clk(cst_30_clk), .rst(cst_30_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_30_in1_valid}), .ready_in_bus({cst_30_in1_ready}), 
		.data_out_bus({cst_30_out1_data}), .valid_out_bus({cst_30_out1_valid}), .ready_out_bus({cst_30_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_86
		(.clk(shl_86_clk), .rst(shl_86_rst),
		.data_in_bus({shl_86_in2_data, shl_86_in1_data}), .valid_in_bus({shl_86_in2_valid, shl_86_in1_valid}), .ready_in_bus({shl_86_in2_ready, shl_86_in1_ready}), 
		.data_out_bus({shl_86_out1_data}), .valid_out_bus({shl_86_out1_valid}), .ready_out_bus({shl_86_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_87
		(.clk(add_87_clk), .rst(add_87_rst),
		.data_in_bus({add_87_in2_data, add_87_in1_data}), .valid_in_bus({add_87_in2_valid, add_87_in1_valid}), .ready_in_bus({add_87_in2_ready, add_87_in1_ready}), 
		.data_out_bus({add_87_out1_data}), .valid_out_bus({add_87_out1_valid}), .ready_out_bus({add_87_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_load_op_load_90
		(.clk(load_90_clk), .rst(load_90_rst),
		.data_in_bus({load_90_in1_data}), .address_in_bus({load_90_in2_data}), .valid_in_bus({load_90_in2_valid, load_90_in1_valid}), .ready_in_bus({load_90_in2_ready, load_90_in1_ready}), 
		.data_out_bus({load_90_out1_data}), .address_out_bus({load_90_out2_data}), .valid_out_bus({load_90_out2_valid, load_90_out1_valid}), .ready_out_bus({load_90_out2_ready, load_90_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_31
		(.clk(cst_31_clk), .rst(cst_31_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_31_in1_valid}), .ready_in_bus({cst_31_in1_ready}), 
		.data_out_bus({cst_31_out1_data}), .valid_out_bus({cst_31_out1_valid}), .ready_out_bus({cst_31_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(7), .DATA_OUT_SIZE(7)) shl_op_shl_91
		(.clk(shl_91_clk), .rst(shl_91_rst),
		.data_in_bus({shl_91_in2_data, shl_91_in1_data}), .valid_in_bus({shl_91_in2_valid, shl_91_in1_valid}), .ready_in_bus({shl_91_in2_ready, shl_91_in1_ready}), 
		.data_out_bus({shl_91_out1_data}), .valid_out_bus({shl_91_out1_valid}), .ready_out_bus({shl_91_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(8), .DATA_OUT_SIZE(8)) add_op_add_92
		(.clk(add_92_clk), .rst(add_92_rst),
		.data_in_bus({add_92_in2_data, add_92_in1_data}), .valid_in_bus({add_92_in2_valid, add_92_in1_valid}), .ready_in_bus({add_92_in2_ready, add_92_in1_ready}), 
		.data_out_bus({add_92_out1_data}), .valid_out_bus({add_92_out1_valid}), .ready_out_bus({add_92_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(8), .DATA_SIZE(32)) mc_load_op_load_95
		(.clk(load_95_clk), .rst(load_95_rst),
		.data_in_bus({load_95_in1_data}), .address_in_bus({load_95_in2_data}), .valid_in_bus({load_95_in2_valid, load_95_in1_valid}), .ready_in_bus({load_95_in2_ready, load_95_in1_ready}), 
		.data_out_bus({load_95_out1_data}), .address_out_bus({load_95_out2_data}), .valid_out_bus({load_95_out2_valid, load_95_out1_valid}), .ready_out_bus({load_95_out2_ready, load_95_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_32
		(.clk(cst_32_clk), .rst(cst_32_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_32_in1_valid}), .ready_in_bus({cst_32_in1_ready}), 
		.data_out_bus({cst_32_out1_data}), .valid_out_bus({cst_32_out1_valid}), .ready_out_bus({cst_32_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) add_op_add_98
		(.clk(add_98_clk), .rst(add_98_rst),
		.data_in_bus({add_98_in2_data, add_98_in1_data}), .valid_in_bus({add_98_in2_valid, add_98_in1_valid}), .ready_in_bus({add_98_in2_ready, add_98_in1_ready}), 
		.data_out_bus({add_98_out1_data}), .valid_out_bus({add_98_out1_valid}), .ready_out_bus({add_98_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) const_node_cst_33
		(.clk(cst_33_clk), .rst(cst_33_rst),
		.data_in_bus({4'd8}), .valid_in_bus({cst_33_in1_valid}), .ready_in_bus({cst_33_in1_ready}), 
		.data_out_bus({cst_33_out1_data}), .valid_out_bus({cst_33_out1_valid}), .ready_out_bus({cst_33_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_99
		(.clk(icmp_99_clk), .rst(icmp_99_rst),
		.data_in_bus({icmp_99_in2_data, icmp_99_in1_data}), .valid_in_bus({icmp_99_in2_valid, icmp_99_in1_valid}), .ready_in_bus({icmp_99_in2_ready, icmp_99_in1_ready}), 
		.data_out_bus({icmp_99_out1_data}), .valid_out_bus({icmp_99_out1_valid}), .ready_out_bus({icmp_99_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n19
		(.clk(phi_n19_clk), .rst(phi_n19_rst),
		.data_in_bus({phi_n19_in2_data, phi_n19_in1_data}), .valid_in_bus({phi_n19_in2_valid, phi_n19_in1_valid}), .ready_in_bus({phi_n19_in2_ready, phi_n19_in1_ready}), 
		.data_out_bus({phi_n19_out1_data}), .valid_out_bus({phi_n19_out1_valid}), .ready_out_bus({phi_n19_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) merge_node_phi_n20
		(.clk(phi_n20_clk), .rst(phi_n20_rst),
		.data_in_bus({phi_n20_in2_data, phi_n20_in1_data}), .valid_in_bus({phi_n20_in2_valid, phi_n20_in1_valid}), .ready_in_bus({phi_n20_in2_ready, phi_n20_in1_ready}), 
		.data_out_bus({phi_n20_out1_data}), .valid_out_bus({phi_n20_out1_valid}), .ready_out_bus({phi_n20_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_13
		(.clk(fork_13_clk), .rst(fork_13_rst),
		.data_in_bus({fork_13_in1_data}), .valid_in_bus({fork_13_in1_valid}), .ready_in_bus({fork_13_in1_ready}), 
		.data_out_bus({fork_13_out3_data, fork_13_out2_data, fork_13_out1_data}), .valid_out_bus({fork_13_out3_valid, fork_13_out2_valid, fork_13_out1_valid}), .ready_out_bus({fork_13_out3_ready, fork_13_out2_ready, fork_13_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_15
		(.clk(fork_15_clk), .rst(fork_15_rst),
		.data_in_bus({fork_15_in1_data}), .valid_in_bus({fork_15_in1_valid}), .ready_in_bus({fork_15_in1_ready}), 
		.data_out_bus({fork_15_out2_data, fork_15_out1_data}), .valid_out_bus({fork_15_out2_valid, fork_15_out1_valid}), .ready_out_bus({fork_15_out2_ready, fork_15_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_31
		(.clk(fork_31_clk), .rst(fork_31_rst),
		.data_in_bus({fork_31_in1_data}), .valid_in_bus({fork_31_in1_valid}), .ready_in_bus({fork_31_in1_ready}), 
		.data_out_bus({fork_31_out2_data, fork_31_out1_data}), .valid_out_bus({fork_31_out2_valid, fork_31_out1_valid}), .ready_out_bus({fork_31_out2_ready, fork_31_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) fork_node_fork_32
		(.clk(fork_32_clk), .rst(fork_32_rst),
		.data_in_bus({fork_32_in1_data}), .valid_in_bus({fork_32_in1_valid}), .ready_in_bus({fork_32_in1_ready}), 
		.data_out_bus({fork_32_out2_data, fork_32_out1_data}), .valid_out_bus({fork_32_out2_valid, fork_32_out1_valid}), .ready_out_bus({fork_32_out2_ready, fork_32_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_35
		(.clk(branch_35_clk), .rst(branch_35_rst),
		.data_in_bus({{31'b0, branch_35_in2_data}, branch_35_in1_data}), .valid_in_bus({branch_35_in2_valid, branch_35_in1_valid}), .ready_in_bus({branch_35_in2_ready, branch_35_in1_ready}), 
		.data_out_bus({branch_35_out2_data, branch_35_out1_data}), .valid_out_bus({branch_35_out2_valid, branch_35_out1_valid}), .ready_out_bus({branch_35_out2_ready, branch_35_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_36
		(.clk(branch_36_clk), .rst(branch_36_rst),
		.data_in_bus({{3'b0, branch_36_in2_data}, branch_36_in1_data}), .valid_in_bus({branch_36_in2_valid, branch_36_in1_valid}), .ready_in_bus({branch_36_in2_ready, branch_36_in1_ready}), 
		.data_out_bus({branch_36_out2_data, branch_36_out1_data}), .valid_out_bus({branch_36_out2_valid, branch_36_out1_valid}), .ready_out_bus({branch_36_out2_ready, branch_36_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_37
		(.clk(branch_37_clk), .rst(branch_37_rst),
		.data_in_bus({{3'b0, branch_37_in2_data}, branch_37_in1_data}), .valid_in_bus({branch_37_in2_valid, branch_37_in1_valid}), .ready_in_bus({branch_37_in2_ready, branch_37_in1_ready}), 
		.data_out_bus({branch_37_out2_data, branch_37_out1_data}), .valid_out_bus({branch_37_out2_valid, branch_37_out1_valid}), .ready_out_bus({branch_37_out2_ready, branch_37_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_38
		(.clk(branch_38_clk), .rst(branch_38_rst),
		.data_in_bus({{3'b0, branch_38_in2_data}, branch_38_in1_data}), .valid_in_bus({branch_38_in2_valid, branch_38_in1_valid}), .ready_in_bus({branch_38_in2_ready, branch_38_in1_ready}), 
		.data_out_bus({branch_38_out2_data, branch_38_out1_data}), .valid_out_bus({branch_38_out2_valid, branch_38_out1_valid}), .ready_out_bus({branch_38_out2_ready, branch_38_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_48
		(.clk(fork_48_clk), .rst(fork_48_rst),
		.data_in_bus({fork_48_in1_data}), .valid_in_bus({fork_48_in1_valid}), .ready_in_bus({fork_48_in1_ready}), 
		.data_out_bus({fork_48_out5_data, fork_48_out4_data, fork_48_out3_data, fork_48_out2_data, fork_48_out1_data}), .valid_out_bus({fork_48_out5_valid, fork_48_out4_valid, fork_48_out3_valid, fork_48_out2_valid, fork_48_out1_valid}), .ready_out_bus({fork_48_out5_ready, fork_48_out4_ready, fork_48_out3_ready, fork_48_out2_ready, fork_48_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_35
		(.clk(phiC_35_clk), .rst(phiC_35_rst),
		.data_in_bus({phiC_35_in2_data, phiC_35_in1_data}), .valid_in_bus({phiC_35_in2_valid, phiC_35_in1_valid}), .ready_in_bus({phiC_35_in2_ready, phiC_35_in1_ready}), 
		.data_out_bus({phiC_35_out2_data, phiC_35_out1_data}), .valid_out_bus({phiC_35_out2_valid, phiC_35_out1_valid}), .ready_out_bus({phiC_35_out2_ready, phiC_35_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_57
		(.clk(branchC_57_clk), .rst(branchC_57_rst),
		.data_in_bus({{branchC_57_in2_data}, branchC_57_in1_data}), .valid_in_bus({branchC_57_in2_valid, branchC_57_in1_valid}), .ready_in_bus({branchC_57_in2_ready, branchC_57_in1_ready}), 
		.data_out_bus({branchC_57_out2_data, branchC_57_out1_data}), .valid_out_bus({branchC_57_out2_valid, branchC_57_out1_valid}), .ready_out_bus({branchC_57_out2_ready, branchC_57_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_21
		(.clk(source_21_clk), .rst(source_21_rst),
		.data_out_bus({source_21_out1_data}), .valid_out_bus({source_21_out1_valid}), .ready_out_bus({source_21_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_22
		(.clk(source_22_clk), .rst(source_22_rst),
		.data_out_bus({source_22_out1_data}), .valid_out_bus({source_22_out1_valid}), .ready_out_bus({source_22_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_23
		(.clk(source_23_clk), .rst(source_23_rst),
		.data_out_bus({source_23_out1_data}), .valid_out_bus({source_23_out1_valid}), .ready_out_bus({source_23_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(4))source_node_source_24
		(.clk(source_24_clk), .rst(source_24_rst),
		.data_out_bus({source_24_out1_data}), .valid_out_bus({source_24_out1_valid}), .ready_out_bus({source_24_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_85
		(.clk(fork_85_clk), .rst(fork_85_rst),
		.data_in_bus({fork_85_in1_data}), .valid_in_bus({fork_85_in1_valid}), .ready_in_bus({fork_85_in1_ready}), 
		.data_out_bus({fork_85_out2_data, fork_85_out1_data}), .valid_out_bus({fork_85_out2_valid, fork_85_out1_valid}), .ready_out_bus({fork_85_out2_ready, fork_85_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4), .COND_SIZE(1)) mux_node_phi_1
		(.clk(phi_1_clk), .rst(phi_1_rst),
		.data_in_bus({{3'b0, phi_1_in1_data}, phi_1_in3_data, phi_1_in2_data}), .valid_in_bus({phi_1_in1_valid, phi_1_in3_valid, phi_1_in2_valid}), .ready_in_bus({phi_1_in1_ready, phi_1_in3_ready, phi_1_in2_ready}), 
		.data_out_bus({phi_1_out1_data}), .valid_out_bus({phi_1_out1_valid}), .ready_out_bus({phi_1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block2
		(.clk(brCst_block2_clk), .rst(brCst_block2_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block2_in1_valid}), .ready_in_bus({brCst_block2_in1_ready}), 
		.data_out_bus({brCst_block2_out1_data}), .valid_out_bus({brCst_block2_out1_valid}), .ready_out_bus({brCst_block2_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_1
		(.clk(cst_1_clk), .rst(cst_1_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_1_in1_valid}), .ready_in_bus({cst_1_in1_ready}), 
		.data_out_bus({cst_1_out1_data}), .valid_out_bus({cst_1_out1_valid}), .ready_out_bus({cst_1_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_1
		(.clk(branch_1_clk), .rst(branch_1_rst),
		.data_in_bus({{branch_1_in2_data}, branch_1_in1_data}), .valid_in_bus({branch_1_in2_valid, branch_1_in1_valid}), .ready_in_bus({branch_1_in2_ready, branch_1_in1_ready}), 
		.data_out_bus({branch_1_out2_data, branch_1_out1_data}), .valid_out_bus({branch_1_out2_valid, branch_1_out1_valid}), .ready_out_bus({branch_1_out2_ready, branch_1_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(4), .DATA_OUT_SIZE(4)) branch_node_branch_2
		(.clk(branch_2_clk), .rst(branch_2_rst),
		.data_in_bus({{3'b0, branch_2_in2_data}, branch_2_in1_data}), .valid_in_bus({branch_2_in2_valid, branch_2_in1_valid}), .ready_in_bus({branch_2_in2_ready, branch_2_in1_ready}), 
		.data_out_bus({branch_2_out2_data, branch_2_out1_data}), .valid_out_bus({branch_2_out2_valid, branch_2_out1_valid}), .ready_out_bus({branch_2_out2_ready, branch_2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_34
		(.clk(fork_34_clk), .rst(fork_34_rst),
		.data_in_bus({fork_34_in1_data}), .valid_in_bus({fork_34_in1_valid}), .ready_in_bus({fork_34_in1_ready}), 
		.data_out_bus({fork_34_out3_data, fork_34_out2_data, fork_34_out1_data}), .valid_out_bus({fork_34_out3_valid, fork_34_out2_valid, fork_34_out1_valid}), .ready_out_bus({fork_34_out3_ready, fork_34_out2_ready, fork_34_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_21
		(.clk(phiC_21_clk), .rst(phiC_21_rst),
		.data_in_bus({phiC_21_in2_data, phiC_21_in1_data}), .valid_in_bus({phiC_21_in2_valid, phiC_21_in1_valid}), .ready_in_bus({phiC_21_in2_ready, phiC_21_in1_ready}), 
		.data_out_bus({phiC_21_out2_data, phiC_21_out1_data}), .valid_out_bus({phiC_21_out2_valid, phiC_21_out1_valid}), .ready_out_bus({phiC_21_out2_ready, phiC_21_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_54
		(.clk(forkC_54_clk), .rst(forkC_54_rst),
		.data_in_bus({forkC_54_in1_data}), .valid_in_bus({forkC_54_in1_valid}), .ready_in_bus({forkC_54_in1_ready}), 
		.data_out_bus({forkC_54_out3_data, forkC_54_out2_data, forkC_54_out1_data}), .valid_out_bus({forkC_54_out3_valid, forkC_54_out2_valid, forkC_54_out1_valid}), .ready_out_bus({forkC_54_out3_ready, forkC_54_out2_ready, forkC_54_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_43
		(.clk(branchC_43_clk), .rst(branchC_43_rst),
		.data_in_bus({{branchC_43_in2_data}, branchC_43_in1_data}), .valid_in_bus({branchC_43_in2_valid, branchC_43_in1_valid}), .ready_in_bus({branchC_43_in2_ready, branchC_43_in1_ready}), 
		.data_out_bus({branchC_43_out2_data, branchC_43_out1_data}), .valid_out_bus({branchC_43_out2_valid, branchC_43_out1_valid}), .ready_out_bus({branchC_43_out2_ready, branchC_43_out1_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(8), .BB_COUNT(1), .LOAD_COUNT(2), .STORE_COUNT(1))MemCont_MC_E
		(.clk(MC_E_clk), .rst(MC_E_rst),
		.io_storeDataOut(E_dout0), .io_storeAddrOut(E_address0), .io_storeEnable(E_we0),
		.io_loadDataIn(E_din1), .io_loadAddrOut(E_address1), .io_loadEnable(E_ce1),
		.io_bbpValids({MC_E_in1_valid}), .io_bb_stCountArray({MC_E_in1_data}), .io_bbReadyToPrevs({MC_E_in1_ready}), .io_rdPortsPrev_ready({MC_E_in5_ready, MC_E_in2_ready}), .io_rdPortsPrev_valid({MC_E_in5_valid, MC_E_in2_valid}), .io_rdPortsPrev_bits({MC_E_in5_data, MC_E_in2_data}), 	
	.io_wrAddrPorts_ready({MC_E_in3_ready}), .io_wrAddrPorts_valid({MC_E_in3_valid}), .io_wrAddrPorts_bits({MC_E_in3_data}), 	
	.io_wrDataPorts_ready({MC_E_in4_ready}), .io_wrDataPorts_valid({MC_E_in4_valid}), .io_wrDataPorts_bits({MC_E_in4_data}), 	
	.io_rdPortsNext_ready({MC_E_out2_ready, MC_E_out1_ready}), .io_rdPortsNext_valid({MC_E_out2_valid, MC_E_out1_valid}), .io_rdPortsNext_bits({MC_E_out2_data, MC_E_out1_data}), 	
	.io_Empty_Valid({MC_E_out3_valid}), .io_Empty_Ready({MC_E_out3_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(8), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_A
		(.clk(MC_A_clk), .rst(MC_A_rst),
		.io_storeDataOut(A_dout0), .io_storeAddrOut(A_address0), .io_storeEnable(A_we0),
		.io_loadDataIn(A_din1), .io_loadAddrOut(A_address1), .io_loadEnable(A_ce1),
		.io_bbpValids({MC_A_in2_valid}), .io_bb_stCountArray({MC_A_in2_data}), .io_bbReadyToPrevs({MC_A_in2_ready}), .io_rdPortsPrev_ready({MC_A_in1_ready}), .io_rdPortsPrev_valid({MC_A_in1_valid}), .io_rdPortsPrev_bits({MC_A_in1_data}), 	
	.io_wrAddrPorts_ready({MC_A_in3_ready}), .io_wrAddrPorts_valid({MC_A_in3_valid}), .io_wrAddrPorts_bits({MC_A_in3_data}), 	
	.io_wrDataPorts_ready({MC_A_in4_ready}), .io_wrDataPorts_valid({MC_A_in4_valid}), .io_wrDataPorts_bits({MC_A_in4_data}), 	
	.io_rdPortsNext_ready({MC_A_out1_ready}), .io_rdPortsNext_valid({MC_A_out1_valid}), .io_rdPortsNext_bits({MC_A_out1_data}), 	
	.io_Empty_Valid({MC_A_out2_valid}), .io_Empty_Ready({MC_A_out2_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(8), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_B
		(.clk(MC_B_clk), .rst(MC_B_rst),
		.io_storeDataOut(B_dout0), .io_storeAddrOut(B_address0), .io_storeEnable(B_we0),
		.io_loadDataIn(B_din1), .io_loadAddrOut(B_address1), .io_loadEnable(B_ce1),
		.io_bbpValids({MC_B_in2_valid}), .io_bb_stCountArray({MC_B_in2_data}), .io_bbReadyToPrevs({MC_B_in2_ready}), .io_rdPortsPrev_ready({MC_B_in1_ready}), .io_rdPortsPrev_valid({MC_B_in1_valid}), .io_rdPortsPrev_bits({MC_B_in1_data}), 	
	.io_wrAddrPorts_ready({MC_B_in3_ready}), .io_wrAddrPorts_valid({MC_B_in3_valid}), .io_wrAddrPorts_bits({MC_B_in3_data}), 	
	.io_wrDataPorts_ready({MC_B_in4_ready}), .io_wrDataPorts_valid({MC_B_in4_valid}), .io_wrDataPorts_bits({MC_B_in4_data}), 	
	.io_rdPortsNext_ready({MC_B_out1_ready}), .io_rdPortsNext_valid({MC_B_out1_valid}), .io_rdPortsNext_bits({MC_B_out1_data}), 	
	.io_Empty_Valid({MC_B_out2_valid}), .io_Empty_Ready({MC_B_out2_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(8), .BB_COUNT(1), .LOAD_COUNT(2), .STORE_COUNT(1))MemCont_MC_F
		(.clk(MC_F_clk), .rst(MC_F_rst),
		.io_storeDataOut(F_dout0), .io_storeAddrOut(F_address0), .io_storeEnable(F_we0),
		.io_loadDataIn(F_din1), .io_loadAddrOut(F_address1), .io_loadEnable(F_ce1),
		.io_bbpValids({MC_F_in1_valid}), .io_bb_stCountArray({MC_F_in1_data}), .io_bbReadyToPrevs({MC_F_in1_ready}), .io_rdPortsPrev_ready({MC_F_in5_ready, MC_F_in2_ready}), .io_rdPortsPrev_valid({MC_F_in5_valid, MC_F_in2_valid}), .io_rdPortsPrev_bits({MC_F_in5_data, MC_F_in2_data}), 	
	.io_wrAddrPorts_ready({MC_F_in3_ready}), .io_wrAddrPorts_valid({MC_F_in3_valid}), .io_wrAddrPorts_bits({MC_F_in3_data}), 	
	.io_wrDataPorts_ready({MC_F_in4_ready}), .io_wrDataPorts_valid({MC_F_in4_valid}), .io_wrDataPorts_bits({MC_F_in4_data}), 	
	.io_rdPortsNext_ready({MC_F_out2_ready, MC_F_out1_ready}), .io_rdPortsNext_valid({MC_F_out2_valid, MC_F_out1_valid}), .io_rdPortsNext_bits({MC_F_out2_data, MC_F_out1_data}), 	
	.io_Empty_Valid({MC_F_out3_valid}), .io_Empty_Ready({MC_F_out3_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(8), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_C
		(.clk(MC_C_clk), .rst(MC_C_rst),
		.io_storeDataOut(C_dout0), .io_storeAddrOut(C_address0), .io_storeEnable(C_we0),
		.io_loadDataIn(C_din1), .io_loadAddrOut(C_address1), .io_loadEnable(C_ce1),
		.io_bbpValids({MC_C_in2_valid}), .io_bb_stCountArray({MC_C_in2_data}), .io_bbReadyToPrevs({MC_C_in2_ready}), .io_rdPortsPrev_ready({MC_C_in1_ready}), .io_rdPortsPrev_valid({MC_C_in1_valid}), .io_rdPortsPrev_bits({MC_C_in1_data}), 	
	.io_wrAddrPorts_ready({MC_C_in3_ready}), .io_wrAddrPorts_valid({MC_C_in3_valid}), .io_wrAddrPorts_bits({MC_C_in3_data}), 	
	.io_wrDataPorts_ready({MC_C_in4_ready}), .io_wrDataPorts_valid({MC_C_in4_valid}), .io_wrDataPorts_bits({MC_C_in4_data}), 	
	.io_rdPortsNext_ready({MC_C_out1_ready}), .io_rdPortsNext_valid({MC_C_out1_valid}), .io_rdPortsNext_bits({MC_C_out1_data}), 	
	.io_Empty_Valid({MC_C_out2_valid}), .io_Empty_Ready({MC_C_out2_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(8), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_D
		(.clk(MC_D_clk), .rst(MC_D_rst),
		.io_storeDataOut(D_dout0), .io_storeAddrOut(D_address0), .io_storeEnable(D_we0),
		.io_loadDataIn(D_din1), .io_loadAddrOut(D_address1), .io_loadEnable(D_ce1),
		.io_bbpValids({MC_D_in2_valid}), .io_bb_stCountArray({MC_D_in2_data}), .io_bbReadyToPrevs({MC_D_in2_ready}), .io_rdPortsPrev_ready({MC_D_in1_ready}), .io_rdPortsPrev_valid({MC_D_in1_valid}), .io_rdPortsPrev_bits({MC_D_in1_data}), 	
	.io_wrAddrPorts_ready({MC_D_in3_ready}), .io_wrAddrPorts_valid({MC_D_in3_valid}), .io_wrAddrPorts_bits({MC_D_in3_data}), 	
	.io_wrDataPorts_ready({MC_D_in4_ready}), .io_wrDataPorts_valid({MC_D_in4_valid}), .io_wrDataPorts_bits({MC_D_in4_data}), 	
	.io_rdPortsNext_ready({MC_D_out1_ready}), .io_rdPortsNext_valid({MC_D_out1_valid}), .io_rdPortsNext_bits({MC_D_out1_data}), 	
	.io_Empty_Valid({MC_D_out2_valid}), .io_Empty_Ready({MC_D_out2_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(8), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_G
		(.clk(MC_G_clk), .rst(MC_G_rst),
		.io_storeDataOut(G_dout0), .io_storeAddrOut(G_address0), .io_storeEnable(G_we0),
		.io_loadDataIn(G_din1), .io_loadAddrOut(G_address1), .io_loadEnable(G_ce1),
		.io_bbpValids({MC_G_in1_valid}), .io_bb_stCountArray({MC_G_in1_data}), .io_bbReadyToPrevs({MC_G_in1_ready}), .io_rdPortsPrev_ready({MC_G_in2_ready}), .io_rdPortsPrev_valid({MC_G_in2_valid}), .io_rdPortsPrev_bits({MC_G_in2_data}), 	
	.io_wrAddrPorts_ready({MC_G_in3_ready}), .io_wrAddrPorts_valid({MC_G_in3_valid}), .io_wrAddrPorts_bits({MC_G_in3_data}), 	
	.io_wrDataPorts_ready({MC_G_in4_ready}), .io_wrDataPorts_valid({MC_G_in4_valid}), .io_wrDataPorts_bits({MC_G_in4_data}), 	
	.io_rdPortsNext_ready({MC_G_out1_ready}), .io_rdPortsNext_valid({MC_G_out1_valid}), .io_rdPortsNext_bits({MC_G_out1_data}), 	
	.io_Empty_Valid({MC_G_out2_valid}), .io_Empty_Ready({MC_G_out2_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_0
		(.clk(sink_0_clk), .rst(sink_0_rst),
		.data_in_bus({sink_0_in1_data}), .valid_in_bus({sink_0_in1_valid}), .ready_in_bus({sink_0_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_1
		(.clk(sink_1_clk), .rst(sink_1_rst),
		.data_in_bus({sink_1_in1_data}), .valid_in_bus({sink_1_in1_valid}), .ready_in_bus({sink_1_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_2
		(.clk(sink_2_clk), .rst(sink_2_rst),
		.data_in_bus({sink_2_in1_data}), .valid_in_bus({sink_2_in1_valid}), .ready_in_bus({sink_2_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_3
		(.clk(sink_3_clk), .rst(sink_3_rst),
		.data_in_bus({sink_3_in1_data}), .valid_in_bus({sink_3_in1_valid}), .ready_in_bus({sink_3_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_4
		(.clk(sink_4_clk), .rst(sink_4_rst),
		.data_in_bus({sink_4_in1_data}), .valid_in_bus({sink_4_in1_valid}), .ready_in_bus({sink_4_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_5
		(.clk(sink_5_clk), .rst(sink_5_rst),
		.data_in_bus({sink_5_in1_data}), .valid_in_bus({sink_5_in1_valid}), .ready_in_bus({sink_5_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_6
		(.clk(sink_6_clk), .rst(sink_6_rst),
		.data_in_bus({sink_6_in1_data}), .valid_in_bus({sink_6_in1_valid}), .ready_in_bus({sink_6_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_7
		(.clk(sink_7_clk), .rst(sink_7_rst),
		.data_in_bus({sink_7_in1_data}), .valid_in_bus({sink_7_in1_valid}), .ready_in_bus({sink_7_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_8
		(.clk(sink_8_clk), .rst(sink_8_rst),
		.data_in_bus({sink_8_in1_data}), .valid_in_bus({sink_8_in1_valid}), .ready_in_bus({sink_8_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_9
		(.clk(sink_9_clk), .rst(sink_9_rst),
		.data_in_bus({sink_9_in1_data}), .valid_in_bus({sink_9_in1_valid}), .ready_in_bus({sink_9_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_10
		(.clk(sink_10_clk), .rst(sink_10_rst),
		.data_in_bus({sink_10_in1_data}), .valid_in_bus({sink_10_in1_valid}), .ready_in_bus({sink_10_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_11
		(.clk(sink_11_clk), .rst(sink_11_rst),
		.data_in_bus({sink_11_in1_data}), .valid_in_bus({sink_11_in1_valid}), .ready_in_bus({sink_11_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_12
		(.clk(sink_12_clk), .rst(sink_12_rst),
		.data_in_bus({sink_12_in1_data}), .valid_in_bus({sink_12_in1_valid}), .ready_in_bus({sink_12_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_13
		(.clk(sink_13_clk), .rst(sink_13_rst),
		.data_in_bus({sink_13_in1_data}), .valid_in_bus({sink_13_in1_valid}), .ready_in_bus({sink_13_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_14
		(.clk(sink_14_clk), .rst(sink_14_rst),
		.data_in_bus({sink_14_in1_data}), .valid_in_bus({sink_14_in1_valid}), .ready_in_bus({sink_14_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_15
		(.clk(sink_15_clk), .rst(sink_15_rst),
		.data_in_bus({sink_15_in1_data}), .valid_in_bus({sink_15_in1_valid}), .ready_in_bus({sink_15_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_16
		(.clk(sink_16_clk), .rst(sink_16_rst),
		.data_in_bus({sink_16_in1_data}), .valid_in_bus({sink_16_in1_valid}), .ready_in_bus({sink_16_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_17
		(.clk(sink_17_clk), .rst(sink_17_rst),
		.data_in_bus({sink_17_in1_data}), .valid_in_bus({sink_17_in1_valid}), .ready_in_bus({sink_17_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_18
		(.clk(sink_18_clk), .rst(sink_18_rst),
		.data_in_bus({sink_18_in1_data}), .valid_in_bus({sink_18_in1_valid}), .ready_in_bus({sink_18_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_19
		(.clk(sink_19_clk), .rst(sink_19_rst),
		.data_in_bus({sink_19_in1_data}), .valid_in_bus({sink_19_in1_valid}), .ready_in_bus({sink_19_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_20
		(.clk(sink_20_clk), .rst(sink_20_rst),
		.data_in_bus({sink_20_in1_data}), .valid_in_bus({sink_20_in1_valid}), .ready_in_bus({sink_20_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_21
		(.clk(sink_21_clk), .rst(sink_21_rst),
		.data_in_bus({sink_21_in1_data}), .valid_in_bus({sink_21_in1_valid}), .ready_in_bus({sink_21_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_22
		(.clk(sink_22_clk), .rst(sink_22_rst),
		.data_in_bus({sink_22_in1_data}), .valid_in_bus({sink_22_in1_valid}), .ready_in_bus({sink_22_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_23
		(.clk(sink_23_clk), .rst(sink_23_rst),
		.data_in_bus({sink_23_in1_data}), .valid_in_bus({sink_23_in1_valid}), .ready_in_bus({sink_23_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_24
		(.clk(sink_24_clk), .rst(sink_24_rst),
		.data_in_bus({sink_24_in1_data}), .valid_in_bus({sink_24_in1_valid}), .ready_in_bus({sink_24_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_25
		(.clk(sink_25_clk), .rst(sink_25_rst),
		.data_in_bus({sink_25_in1_data}), .valid_in_bus({sink_25_in1_valid}), .ready_in_bus({sink_25_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_26
		(.clk(sink_26_clk), .rst(sink_26_rst),
		.data_in_bus({sink_26_in1_data}), .valid_in_bus({sink_26_in1_valid}), .ready_in_bus({sink_26_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_27
		(.clk(sink_27_clk), .rst(sink_27_rst),
		.data_in_bus({sink_27_in1_data}), .valid_in_bus({sink_27_in1_valid}), .ready_in_bus({sink_27_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_28
		(.clk(sink_28_clk), .rst(sink_28_rst),
		.data_in_bus({sink_28_in1_data}), .valid_in_bus({sink_28_in1_valid}), .ready_in_bus({sink_28_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(4))sink_node_sink_29
		(.clk(sink_29_clk), .rst(sink_29_rst),
		.data_in_bus({sink_29_in1_data}), .valid_in_bus({sink_29_in1_valid}), .ready_in_bus({sink_29_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_30
		(.clk(sink_30_clk), .rst(sink_30_rst),
		.data_in_bus({sink_30_in1_data}), .valid_in_bus({sink_30_in1_valid}), .ready_in_bus({sink_30_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_31
		(.clk(sink_31_clk), .rst(sink_31_rst),
		.data_in_bus({sink_31_in1_data}), .valid_in_bus({sink_31_in1_valid}), .ready_in_bus({sink_31_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_32
		(.clk(sink_32_clk), .rst(sink_32_rst),
		.data_in_bus({sink_32_in1_data}), .valid_in_bus({sink_32_in1_valid}), .ready_in_bus({sink_32_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_33
		(.clk(sink_33_clk), .rst(sink_33_rst),
		.data_in_bus({sink_33_in1_data}), .valid_in_bus({sink_33_in1_valid}), .ready_in_bus({sink_33_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_34
		(.clk(sink_34_clk), .rst(sink_34_rst),
		.data_in_bus({sink_34_in1_data}), .valid_in_bus({sink_34_in1_valid}), .ready_in_bus({sink_34_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_35
		(.clk(sink_35_clk), .rst(sink_35_rst),
		.data_in_bus({sink_35_in1_data}), .valid_in_bus({sink_35_in1_valid}), .ready_in_bus({sink_35_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_36
		(.clk(sink_36_clk), .rst(sink_36_rst),
		.data_in_bus({sink_36_in1_data}), .valid_in_bus({sink_36_in1_valid}), .ready_in_bus({sink_36_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_37
		(.clk(sink_37_clk), .rst(sink_37_rst),
		.data_in_bus({sink_37_in1_data}), .valid_in_bus({sink_37_in1_valid}), .ready_in_bus({sink_37_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_38
		(.clk(sink_38_clk), .rst(sink_38_rst),
		.data_in_bus({sink_38_in1_data}), .valid_in_bus({sink_38_in1_valid}), .ready_in_bus({sink_38_in1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_100
		(.clk(Buffer_100_clk), .rst(Buffer_100_rst),
		.data_in_bus({Buffer_100_in1_data}), .valid_in_bus({Buffer_100_in1_valid}), .ready_in_bus({Buffer_100_in1_ready}), 
		.data_out_bus({Buffer_100_out1_data}), .valid_out_bus({Buffer_100_out1_valid}), .ready_out_bus({Buffer_100_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_101
		(.clk(Buffer_101_clk), .rst(Buffer_101_rst),
		.data_in_bus({Buffer_101_in1_data}), .valid_in_bus({Buffer_101_in1_valid}), .ready_in_bus({Buffer_101_in1_ready}), 
		.data_out_bus({Buffer_101_out1_data}), .valid_out_bus({Buffer_101_out1_valid}), .ready_out_bus({Buffer_101_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_102
		(.clk(Buffer_102_clk), .rst(Buffer_102_rst),
		.data_in_bus({Buffer_102_in1_data}), .valid_in_bus({Buffer_102_in1_valid}), .ready_in_bus({Buffer_102_in1_ready}), 
		.data_out_bus({Buffer_102_out1_data}), .valid_out_bus({Buffer_102_out1_valid}), .ready_out_bus({Buffer_102_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_103
		(.clk(Buffer_103_clk), .rst(Buffer_103_rst),
		.data_in_bus({Buffer_103_in1_data}), .valid_in_bus({Buffer_103_in1_valid}), .ready_in_bus({Buffer_103_in1_ready}), 
		.data_out_bus({Buffer_103_out1_data}), .valid_out_bus({Buffer_103_out1_valid}), .ready_out_bus({Buffer_103_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_104
		(.clk(Buffer_104_clk), .rst(Buffer_104_rst),
		.data_in_bus({Buffer_104_in1_data}), .valid_in_bus({Buffer_104_in1_valid}), .ready_in_bus({Buffer_104_in1_ready}), 
		.data_out_bus({Buffer_104_out1_data}), .valid_out_bus({Buffer_104_out1_valid}), .ready_out_bus({Buffer_104_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_105
		(.clk(Buffer_105_clk), .rst(Buffer_105_rst),
		.data_in_bus({Buffer_105_in1_data}), .valid_in_bus({Buffer_105_in1_valid}), .ready_in_bus({Buffer_105_in1_ready}), 
		.data_out_bus({Buffer_105_out1_data}), .valid_out_bus({Buffer_105_out1_valid}), .ready_out_bus({Buffer_105_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_106
		(.clk(Buffer_106_clk), .rst(Buffer_106_rst),
		.data_in_bus({Buffer_106_in1_data}), .valid_in_bus({Buffer_106_in1_valid}), .ready_in_bus({Buffer_106_in1_ready}), 
		.data_out_bus({Buffer_106_out1_data}), .valid_out_bus({Buffer_106_out1_valid}), .ready_out_bus({Buffer_106_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_107
		(.clk(Buffer_107_clk), .rst(Buffer_107_rst),
		.data_in_bus({Buffer_107_in1_data}), .valid_in_bus({Buffer_107_in1_valid}), .ready_in_bus({Buffer_107_in1_ready}), 
		.data_out_bus({Buffer_107_out1_data}), .valid_out_bus({Buffer_107_out1_valid}), .ready_out_bus({Buffer_107_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_108
		(.clk(Buffer_108_clk), .rst(Buffer_108_rst),
		.data_in_bus({Buffer_108_in1_data}), .valid_in_bus({Buffer_108_in1_valid}), .ready_in_bus({Buffer_108_in1_ready}), 
		.data_out_bus({Buffer_108_out1_data}), .valid_out_bus({Buffer_108_out1_valid}), .ready_out_bus({Buffer_108_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_109
		(.clk(Buffer_109_clk), .rst(Buffer_109_rst),
		.data_in_bus({Buffer_109_in1_data}), .valid_in_bus({Buffer_109_in1_valid}), .ready_in_bus({Buffer_109_in1_ready}), 
		.data_out_bus({Buffer_109_out1_data}), .valid_out_bus({Buffer_109_out1_valid}), .ready_out_bus({Buffer_109_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_110
		(.clk(Buffer_110_clk), .rst(Buffer_110_rst),
		.data_in_bus({Buffer_110_in1_data}), .valid_in_bus({Buffer_110_in1_valid}), .ready_in_bus({Buffer_110_in1_ready}), 
		.data_out_bus({Buffer_110_out1_data}), .valid_out_bus({Buffer_110_out1_valid}), .ready_out_bus({Buffer_110_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_111
		(.clk(Buffer_111_clk), .rst(Buffer_111_rst),
		.data_in_bus({Buffer_111_in1_data}), .valid_in_bus({Buffer_111_in1_valid}), .ready_in_bus({Buffer_111_in1_ready}), 
		.data_out_bus({Buffer_111_out1_data}), .valid_out_bus({Buffer_111_out1_valid}), .ready_out_bus({Buffer_111_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_112
		(.clk(Buffer_112_clk), .rst(Buffer_112_rst),
		.data_in_bus({Buffer_112_in1_data}), .valid_in_bus({Buffer_112_in1_valid}), .ready_in_bus({Buffer_112_in1_ready}), 
		.data_out_bus({Buffer_112_out1_data}), .valid_out_bus({Buffer_112_out1_valid}), .ready_out_bus({Buffer_112_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_113
		(.clk(Buffer_113_clk), .rst(Buffer_113_rst),
		.data_in_bus({Buffer_113_in1_data}), .valid_in_bus({Buffer_113_in1_valid}), .ready_in_bus({Buffer_113_in1_ready}), 
		.data_out_bus({Buffer_113_out1_data}), .valid_out_bus({Buffer_113_out1_valid}), .ready_out_bus({Buffer_113_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_114
		(.clk(Buffer_114_clk), .rst(Buffer_114_rst),
		.data_in_bus({Buffer_114_in1_data}), .valid_in_bus({Buffer_114_in1_valid}), .ready_in_bus({Buffer_114_in1_ready}), 
		.data_out_bus({Buffer_114_out1_data}), .valid_out_bus({Buffer_114_out1_valid}), .ready_out_bus({Buffer_114_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_115
		(.clk(Buffer_115_clk), .rst(Buffer_115_rst),
		.data_in_bus({Buffer_115_in1_data}), .valid_in_bus({Buffer_115_in1_valid}), .ready_in_bus({Buffer_115_in1_ready}), 
		.data_out_bus({Buffer_115_out1_data}), .valid_out_bus({Buffer_115_out1_valid}), .ready_out_bus({Buffer_115_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_116
		(.clk(Buffer_116_clk), .rst(Buffer_116_rst),
		.data_in_bus({Buffer_116_in1_data}), .valid_in_bus({Buffer_116_in1_valid}), .ready_in_bus({Buffer_116_in1_ready}), 
		.data_out_bus({Buffer_116_out1_data}), .valid_out_bus({Buffer_116_out1_valid}), .ready_out_bus({Buffer_116_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_117
		(.clk(Buffer_117_clk), .rst(Buffer_117_rst),
		.data_in_bus({Buffer_117_in1_data}), .valid_in_bus({Buffer_117_in1_valid}), .ready_in_bus({Buffer_117_in1_ready}), 
		.data_out_bus({Buffer_117_out1_data}), .valid_out_bus({Buffer_117_out1_valid}), .ready_out_bus({Buffer_117_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_118
		(.clk(Buffer_118_clk), .rst(Buffer_118_rst),
		.data_in_bus({Buffer_118_in1_data}), .valid_in_bus({Buffer_118_in1_valid}), .ready_in_bus({Buffer_118_in1_ready}), 
		.data_out_bus({Buffer_118_out1_data}), .valid_out_bus({Buffer_118_out1_valid}), .ready_out_bus({Buffer_118_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_119
		(.clk(Buffer_119_clk), .rst(Buffer_119_rst),
		.data_in_bus({Buffer_119_in1_data}), .valid_in_bus({Buffer_119_in1_valid}), .ready_in_bus({Buffer_119_in1_ready}), 
		.data_out_bus({Buffer_119_out1_data}), .valid_out_bus({Buffer_119_out1_valid}), .ready_out_bus({Buffer_119_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_120
		(.clk(Buffer_120_clk), .rst(Buffer_120_rst),
		.data_in_bus({Buffer_120_in1_data}), .valid_in_bus({Buffer_120_in1_valid}), .ready_in_bus({Buffer_120_in1_ready}), 
		.data_out_bus({Buffer_120_out1_data}), .valid_out_bus({Buffer_120_out1_valid}), .ready_out_bus({Buffer_120_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_121
		(.clk(Buffer_121_clk), .rst(Buffer_121_rst),
		.data_in_bus({Buffer_121_in1_data}), .valid_in_bus({Buffer_121_in1_valid}), .ready_in_bus({Buffer_121_in1_ready}), 
		.data_out_bus({Buffer_121_out1_data}), .valid_out_bus({Buffer_121_out1_valid}), .ready_out_bus({Buffer_121_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_122
		(.clk(Buffer_122_clk), .rst(Buffer_122_rst),
		.data_in_bus({Buffer_122_in1_data}), .valid_in_bus({Buffer_122_in1_valid}), .ready_in_bus({Buffer_122_in1_ready}), 
		.data_out_bus({Buffer_122_out1_data}), .valid_out_bus({Buffer_122_out1_valid}), .ready_out_bus({Buffer_122_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_123
		(.clk(Buffer_123_clk), .rst(Buffer_123_rst),
		.data_in_bus({Buffer_123_in1_data}), .valid_in_bus({Buffer_123_in1_valid}), .ready_in_bus({Buffer_123_in1_ready}), 
		.data_out_bus({Buffer_123_out1_data}), .valid_out_bus({Buffer_123_out1_valid}), .ready_out_bus({Buffer_123_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_124
		(.clk(Buffer_124_clk), .rst(Buffer_124_rst),
		.data_in_bus({Buffer_124_in1_data}), .valid_in_bus({Buffer_124_in1_valid}), .ready_in_bus({Buffer_124_in1_ready}), 
		.data_out_bus({Buffer_124_out1_data}), .valid_out_bus({Buffer_124_out1_valid}), .ready_out_bus({Buffer_124_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_125
		(.clk(Buffer_125_clk), .rst(Buffer_125_rst),
		.data_in_bus({Buffer_125_in1_data}), .valid_in_bus({Buffer_125_in1_valid}), .ready_in_bus({Buffer_125_in1_ready}), 
		.data_out_bus({Buffer_125_out1_data}), .valid_out_bus({Buffer_125_out1_valid}), .ready_out_bus({Buffer_125_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_126
		(.clk(Buffer_126_clk), .rst(Buffer_126_rst),
		.data_in_bus({Buffer_126_in1_data}), .valid_in_bus({Buffer_126_in1_valid}), .ready_in_bus({Buffer_126_in1_ready}), 
		.data_out_bus({Buffer_126_out1_data}), .valid_out_bus({Buffer_126_out1_valid}), .ready_out_bus({Buffer_126_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_127
		(.clk(Buffer_127_clk), .rst(Buffer_127_rst),
		.data_in_bus({Buffer_127_in1_data}), .valid_in_bus({Buffer_127_in1_valid}), .ready_in_bus({Buffer_127_in1_ready}), 
		.data_out_bus({Buffer_127_out1_data}), .valid_out_bus({Buffer_127_out1_valid}), .ready_out_bus({Buffer_127_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_128
		(.clk(Buffer_128_clk), .rst(Buffer_128_rst),
		.data_in_bus({Buffer_128_in1_data}), .valid_in_bus({Buffer_128_in1_valid}), .ready_in_bus({Buffer_128_in1_ready}), 
		.data_out_bus({Buffer_128_out1_data}), .valid_out_bus({Buffer_128_out1_valid}), .ready_out_bus({Buffer_128_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_129
		(.clk(Buffer_129_clk), .rst(Buffer_129_rst),
		.data_in_bus({Buffer_129_in1_data}), .valid_in_bus({Buffer_129_in1_valid}), .ready_in_bus({Buffer_129_in1_ready}), 
		.data_out_bus({Buffer_129_out1_data}), .valid_out_bus({Buffer_129_out1_valid}), .ready_out_bus({Buffer_129_out1_ready}));

	and_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) and_op_and_300
		(.clk(and_300_clk), .rst(and_300_rst),
		.data_in_bus({and_300_in2_data, and_300_in1_data}), .valid_in_bus({and_300_in2_valid, and_300_in1_valid}), .ready_in_bus({and_300_in2_ready, and_300_in1_ready}), 
		.data_out_bus({and_300_out1_data}), .valid_out_bus({and_300_out1_valid}), .ready_out_bus({and_300_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_300
		(.clk(Buffer_300_clk), .rst(Buffer_300_rst),
		.data_in_bus({Buffer_300_in1_data}), .valid_in_bus({Buffer_300_in1_valid}), .ready_in_bus({Buffer_300_in1_ready}), 
		.data_out_bus({Buffer_300_out1_data}), .valid_out_bus({Buffer_300_out1_valid}), .ready_out_bus({Buffer_300_out1_ready}));

	and_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) and_op_and_301
		(.clk(and_301_clk), .rst(and_301_rst),
		.data_in_bus({and_301_in2_data, and_301_in1_data}), .valid_in_bus({and_301_in2_valid, and_301_in1_valid}), .ready_in_bus({and_301_in2_ready, and_301_in1_ready}), 
		.data_out_bus({and_301_out1_data}), .valid_out_bus({and_301_out1_valid}), .ready_out_bus({and_301_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_301
		(.clk(Buffer_301_clk), .rst(Buffer_301_rst),
		.data_in_bus({Buffer_301_in1_data}), .valid_in_bus({Buffer_301_in1_valid}), .ready_in_bus({Buffer_301_in1_ready}), 
		.data_out_bus({Buffer_301_out1_data}), .valid_out_bus({Buffer_301_out1_valid}), .ready_out_bus({Buffer_301_out1_ready}));

	and_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) and_op_and_302
		(.clk(and_302_clk), .rst(and_302_rst),
		.data_in_bus({and_302_in2_data, and_302_in1_data}), .valid_in_bus({and_302_in2_valid, and_302_in1_valid}), .ready_in_bus({and_302_in2_ready, and_302_in1_ready}), 
		.data_out_bus({and_302_out1_data}), .valid_out_bus({and_302_out1_valid}), .ready_out_bus({and_302_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_302
		(.clk(Buffer_302_clk), .rst(Buffer_302_rst),
		.data_in_bus({Buffer_302_in1_data}), .valid_in_bus({Buffer_302_in1_valid}), .ready_in_bus({Buffer_302_in1_ready}), 
		.data_out_bus({Buffer_302_out1_data}), .valid_out_bus({Buffer_302_out1_valid}), .ready_out_bus({Buffer_302_out1_ready}));

	and_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) and_op_and_303
		(.clk(and_303_clk), .rst(and_303_rst),
		.data_in_bus({and_303_in2_data, and_303_in1_data}), .valid_in_bus({and_303_in2_valid, and_303_in1_valid}), .ready_in_bus({and_303_in2_ready, and_303_in1_ready}), 
		.data_out_bus({and_303_out1_data}), .valid_out_bus({and_303_out1_valid}), .ready_out_bus({and_303_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_303
		(.clk(Buffer_303_clk), .rst(Buffer_303_rst),
		.data_in_bus({Buffer_303_in1_data}), .valid_in_bus({Buffer_303_in1_valid}), .ready_in_bus({Buffer_303_in1_ready}), 
		.data_out_bus({Buffer_303_out1_data}), .valid_out_bus({Buffer_303_out1_valid}), .ready_out_bus({Buffer_303_out1_ready}));

	and_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) and_op_and_304
		(.clk(and_304_clk), .rst(and_304_rst),
		.data_in_bus({and_304_in2_data, and_304_in1_data}), .valid_in_bus({and_304_in2_valid, and_304_in1_valid}), .ready_in_bus({and_304_in2_ready, and_304_in1_ready}), 
		.data_out_bus({and_304_out1_data}), .valid_out_bus({and_304_out1_valid}), .ready_out_bus({and_304_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_304
		(.clk(Buffer_304_clk), .rst(Buffer_304_rst),
		.data_in_bus({Buffer_304_in1_data}), .valid_in_bus({Buffer_304_in1_valid}), .ready_in_bus({Buffer_304_in1_ready}), 
		.data_out_bus({Buffer_304_out1_data}), .valid_out_bus({Buffer_304_out1_valid}), .ready_out_bus({Buffer_304_out1_ready}));

	and_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) and_op_and_305
		(.clk(and_305_clk), .rst(and_305_rst),
		.data_in_bus({and_305_in2_data, and_305_in1_data}), .valid_in_bus({and_305_in2_valid, and_305_in1_valid}), .ready_in_bus({and_305_in2_ready, and_305_in1_ready}), 
		.data_out_bus({and_305_out1_data}), .valid_out_bus({and_305_out1_valid}), .ready_out_bus({and_305_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_305
		(.clk(Buffer_305_clk), .rst(Buffer_305_rst),
		.data_in_bus({Buffer_305_in1_data}), .valid_in_bus({Buffer_305_in1_valid}), .ready_in_bus({Buffer_305_in1_ready}), 
		.data_out_bus({Buffer_305_out1_data}), .valid_out_bus({Buffer_305_out1_valid}), .ready_out_bus({Buffer_305_out1_ready}));

endmodule

