module gemver(
	input [5 : 0] fork_14__icmp_101__data__0__anchor__in,
	input start_0__forkC_44__ready__0__anchor__in,
	input [5 : 0] fork_4__load_51__data__0__anchor__in,
	input fork_4__add_54__valid__0__anchor__in,
	input [31 : 0] Buffer_23__phi_n27__data__0__anchor__in,
	input branch_7__Buffer_25__valid__0__anchor__in,
	input [31 : 0] load_92__mul_93__data__0__anchor__in,
	input [31 : 0] store_3__MC_w__data__0__anchor__in,
	input branch_43__Buffer_23__ready__0__anchor__in,
	input load_66__MC_x__valid__0__anchor__in,
	input fork_14__branch_45__valid__0__anchor__in,
	input [31 : 0] branch_33__phi_n21__data__0__anchor__in,
	input [31 : 0] z_din1,
	input beta_valid_in,
	input phiC_32__forkC_49__valid__0__anchor__in,
	input load_69__add_70__valid__0__anchor__in,
	input fork_40__branch_37__ready__0__anchor__in,
	input brCst_block2__fork_30__data__0__anchor__in,
	input fork_41__branch_43__valid__0__anchor__in,
	input forkC_51__cst_26__valid__0__anchor__in,
	input [5 : 0] cst_6__add_32__data__0__anchor__in,
	input branchC_52__phiC_34__data__0__anchor__in,
	input [31 : 0] fork_23__mul_48__data__0__anchor__in,
	input [31 : 0] branch_36__sink_25__data__0__anchor__in,
	input branch_0__phi_1__valid__0__anchor__in,
	input phi_n6__branch_9__ready__0__anchor__in,
	input fork_30__branch_5__ready__0__anchor__in,
	input source_4__cst_6__ready__0__anchor__in,
	input Buffer_6__phiC_38__data__0__anchor__in,
	input Buffer_27__phiC_32__valid__0__anchor__in,
	input store_3__MC_w__ready__1__anchor__in,
	input cst_2__shl_4__ready__0__anchor__in,
	input [31 : 0] branch_5__phi_n6__data__0__anchor__in,
	input branch_44__sink_30__ready__0__anchor__in,
	input add_59__fork_7__valid__0__anchor__in,
	input [31 : 0] phi_n19__branch_31__data__0__anchor__in,
	input forkC_45__branchC_47__valid__0__anchor__in,
	input source_4__cst_6__data__0__anchor__in,
	input [31 : 0] branch_5__sink_5__data__0__anchor__in,
	input [31 : 0] store_1__MC_x__data__0__anchor__in,
	input fork_36__branch_29__ready__0__anchor__in,
	input forkC_55__branchC_57__ready__0__anchor__in,
	input fork_17__shl_25__ready__0__anchor__in,
	input branch_5__sink_5__valid__0__anchor__in,
	input branch_29__Buffer_24__valid__0__anchor__in,
	input cst_15__branch_30__data__0__anchor__in,
	input [11 : 0] load_88__MC_A__data__0__anchor__in,
	input [5 : 0] branch_4__phi_n5__data__0__anchor__in,
	input add_29__fork_1__valid__0__anchor__in,
	input fork_40__branch_38__data__0__anchor__in,
	input phi_n11__branch_20__ready__0__anchor__in,
	input branch_3__sink_3__valid__0__anchor__in,
	input mul_15__add_16__ready__0__anchor__in,
	input [5 : 0] load_92__MC_x__data__0__anchor__in,
	input Buffer_12__phi_41__valid__0__anchor__in,
	input MC_z__load_69__ready__0__anchor__in,
	input [5 : 0] fork_8__add_73__data__0__anchor__in,
	input fork_11__load_92__valid__0__anchor__in,
	input Buffer_7__phiC_36__data__0__anchor__in,
	input phiC_34__forkC_51__data__0__anchor__in,
	input [5 : 0] branch_8__phi_n2__data__0__anchor__in,
	input MC_v2__load_22__valid__0__anchor__in,
	input [5 : 0] branch_32__Buffer_10__data__0__anchor__in,
	input fork_40__branch_36__ready__0__anchor__in,
	input forkC_53__branchC_55__ready__0__anchor__in,
	input phi_n23__store_3__ready__0__anchor__in,
	input [31 : 0] u1_din1,
	input phiC_32__forkC_49__data__0__anchor__in,
	input forkC_45__cst_1__ready__0__anchor__in,
	input branch_1__sink_1__ready__0__anchor__in,
	input cst_14__icmp_60__valid__0__anchor__in,
	input [31 : 0] y_din0,
	input Buffer_30__forkC_55__ready__0__anchor__in,
	input phiC_35__forkC_52__valid__0__anchor__in,
	input fork_42__branch_45__data__0__anchor__in,
	input [31 : 0] fork_28__branch_43__data__0__anchor__in,
	input branch_32__Buffer_10__valid__0__anchor__in,
	input fork_38__branchC_55__ready__0__anchor__in,
	input fork_40__branch_39__data__0__anchor__in,
	input [31 : 0] mul_48__mul_52__data__0__anchor__in,
	input branch_31__phi_n20__ready__0__anchor__in,
	input [31 : 0] load_80__branch_36__data__0__anchor__in,
	input [31 : 0] phi_n17__fork_23__data__0__anchor__in,
	input MC_u2__load_19__ready__0__anchor__in,
	input fork_11__add_95__valid__0__anchor__in,
	input fork_38__branch_32__valid__0__anchor__in,
	input fork_23__mul_48__valid__0__anchor__in,
	input forkC_48__brCst_block5__valid__0__anchor__in,
	input MC_u1__load_11__valid__0__anchor__in,
	input phi_n20__branch_33__ready__0__anchor__in,
	input Buffer_24__phi_n11__valid__0__anchor__in,
	input fork_36__branchC_53__valid__0__anchor__in,
	input branchC_59__phiC_41__valid__0__anchor__in,
	input cst_24__icmp_101__valid__0__anchor__in,
	input phiC_36__phi_63__data__0__anchor__in,
	input fork_65__phi_82__data__0__anchor__in,
	input fork_34__branch_17__ready__0__anchor__in,
	input fork_32__branch_11__ready__0__anchor__in,
	input branch_18__sink_13__valid__0__anchor__in,
	input [31 : 0] Buffer_4__phi_n6__data__0__anchor__in,
	input [5 : 0] Buffer_29__phi_83__data__0__anchor__in,
	input fork_38__branch_33__data__0__anchor__in,
	input branch_3__phi_3__ready__0__anchor__in,
	input branch_21__sink_16__valid__0__anchor__in,
	input load_19__mul_23__valid__0__anchor__in,
	input store_3__MC_w__ready__0__anchor__in,
	input [31 : 0] beta__branch_1__data__0__anchor__in,
	input cst_9__branch_18__ready__0__anchor__in,
	input mul_48__mul_52__ready__0__anchor__in,
	input branch_6__phi_n7__ready__0__anchor__in,
	input store_1__MC_x__ready__0__anchor__in,
	input fork_31__branch_9__data__0__anchor__in,
	input [31 : 0] branch_6__sink_6__data__0__anchor__in,
	input fork_38__branchC_55__valid__0__anchor__in,
	input MC_x__end_0__valid__0__anchor__in,
	input [11 : 0] fork_22__add_44__data__0__anchor__in,
	input branch_28__sink_19__valid__0__anchor__in,
	input [11 : 0] load_47__MC_A__data__0__anchor__in,
	input [31 : 0] mul_89__mul_93__data__0__anchor__in,
	input source_3__cst_5__valid__0__anchor__in,
	input brCst_block1__fork_29__data__0__anchor__in,
	input Buffer_6__phiC_38__ready__0__anchor__in,
	input branchC_53__phiC_35__ready__0__anchor__in,
	input branchC_53__phiC_35__valid__0__anchor__in,
	input brCst_block5__fork_33__valid__0__anchor__in,
	input branch_4__sink_4__valid__0__anchor__in,
	input branch_26__Buffer_18__valid__0__anchor__in,
	input branchC_47__phiC_29__data__0__anchor__in,
	input store_2__MC_x__ready__0__anchor__in,
	input fork_0__load_14__valid__0__anchor__in,
	input fork_10__branch_39__ready__0__anchor__in,
	input add_5__load_8__ready__0__anchor__in,
	input [5 : 0] fork_11__load_92__data__0__anchor__in,
	input phiC_32__forkC_49__ready__0__anchor__in,
	input fork_28__branch_43__ready__0__anchor__in,
	input Buffer_2__phiC_39__ready__0__anchor__in,
	input cst_21__add_95__ready__0__anchor__in,
	input [31 : 0] phi_n10__branch_19__data__0__anchor__in,
	input fork_37__branch_30__valid__0__anchor__in,
	input branch_33__phi_n21__valid__0__anchor__in,
	input fork_39__branch_35__data__0__anchor__in,
	input branchC_47__phiC_29__ready__0__anchor__in,
	input add_16__add_24__valid__0__anchor__in,
	input branch_13__phi_n9__valid__0__anchor__in,
	input fork_3__load_39__valid__0__anchor__in,
	input [31 : 0] branch_44__sink_30__data__0__anchor__in,
	input branch_7__Buffer_25__ready__0__anchor__in,
	input forkC_52__brCst_block9__data__0__anchor__in,
	input Buffer_3__phi_42__valid__0__anchor__in,
	input brCst_block5__fork_33__ready__0__anchor__in,
	input [5 : 0] fork_13__icmp_96__data__0__anchor__in,
	input fork_30__branch_6__ready__0__anchor__in,
	input forkC_54__branchC_56__ready__0__anchor__in,
	input cst_23__add_100__ready__0__anchor__in,
	input [31 : 0] branch_26__Buffer_18__data__0__anchor__in,
	input forkC_51__branchC_53__data__0__anchor__in,
	input icmp_60__fork_36__valid__0__anchor__in,
	input load_8__MC_A__valid__0__anchor__in,
	input branch_21__sink_16__ready__0__anchor__in,
	input fork_37__branch_31__valid__0__anchor__in,
	input fork_0__add_29__valid__0__anchor__in,
	input fork_23__mul_48__ready__0__anchor__in,
	input branch_31__sink_21__valid__0__anchor__in,
	input MC_x__load_66__ready__0__anchor__in,
	input source_6__cst_10__ready__0__anchor__in,
	input [5 : 0] fork_2__branch_11__data__0__anchor__in,
	input branch_11__Buffer_26__ready__0__anchor__in,
	input [31 : 0] MC_A__load_47__data__0__anchor__in,
	input fork_13__icmp_96__ready__0__anchor__in,
	input fork_0__add_26__valid__0__anchor__in,
	input [5 : 0] fork_22__branch_24__data__0__anchor__in,
	input fork_37__branch_31__data__0__anchor__in,
	input forkC_45__branchC_47__data__0__anchor__in,
	input branch_18__phi_42__valid__0__anchor__in,
	input fork_17__load_11__ready__0__anchor__in,
	input store_3__MC_w__valid__0__anchor__in,
	input [31 : 0] mul_93__add_94__data__0__anchor__in,
	input fork_7__icmp_60__ready__0__anchor__in,
	input store_0__MC_A__ready__1__anchor__in,
	input [31 : 0] v1_din0,
	input fork_34__branch_18__ready__0__anchor__in,
	input fork_40__branch_37__data__0__anchor__in,
	input fork_40__branch_39__ready__0__anchor__in,
	input store_2__MC_x__valid__0__anchor__in,
	input Buffer_24__phi_n11__ready__0__anchor__in,
	input fork_35__branchC_52__ready__0__anchor__in,
	input source_17__cst_24__valid__0__anchor__in,
	input [5 : 0] source_12__cst_17__data__0__anchor__in,
	input [31 : 0] Buffer_24__phi_n11__data__0__anchor__in,
	input phiC_36__phi_63__ready__0__anchor__in,
	input [31 : 0] x_din1,
	input branch_40__Buffer_8__ready__0__anchor__in,
	input fork_23__branch_25__valid__0__anchor__in,
	input MC_A__end_0__ready__0__anchor__in,
	input load_39__MC_x__valid__0__anchor__in,
	input load_39__MC_x__ready__0__anchor__in,
	input MC_v1__load_14__ready__0__anchor__in,
	input phiC_38__phi_77__ready__0__anchor__in,
	input branch_26__Buffer_18__ready__0__anchor__in,
	input start_in,
	input [2 : 0] source_1__cst_3__data__0__anchor__in,
	input phiC_36__forkC_53__data__0__anchor__in,
	input fork_26__store_3__ready__0__anchor__in,
	input forkC_57__branchC_59__ready__0__anchor__in,
	input branch_9__Buffer_4__ready__0__anchor__in,
	input [31 : 0] branch_31__phi_n20__data__0__anchor__in,
	input [5 : 0] Buffer_10__phi_63__data__0__anchor__in,
	input branch_13__Buffer_19__valid__0__anchor__in,
	input [31 : 0] branch_27__Buffer_13__data__0__anchor__in,
	input [5 : 0] Buffer_14__phi_n5__data__0__anchor__in,
	input cst_20__shl_84__ready__0__anchor__in,
	input branchC_46__phiC_28__ready__0__anchor__in,
	input fork_7__branch_28__ready__0__anchor__in,
	input branchC_59__Buffer_6__ready__0__anchor__in,
	input cst_22__icmp_96__ready__0__anchor__in,
	input fork_65__phi_83__ready__0__anchor__in,
	input branch_9__phi_n3__ready__0__anchor__in,
	input icmp_101__fork_42__ready__0__anchor__in,
	input load_69__MC_z__valid__0__anchor__in,
	input branch_16__sink_11__ready__0__anchor__in,
	input fork_6__icmp_55__ready__0__anchor__in,
	input fork_34__branch_21__ready__0__anchor__in,
	input branchC_47__phiC_29__valid__0__anchor__in,
	input fork_17__branch_8__valid__0__anchor__in,
	input fork_35__branch_25__data__0__anchor__in,
	input forkC_44__cst_0__ready__0__anchor__in,
	input clk,
	input fork_35__branchC_52__data__0__anchor__in,
	input branch_26__phi_n15__valid__0__anchor__in,
	input [31 : 0] phi_n9__branch_16__data__0__anchor__in,
	input [31 : 0] phi_n18__branch_26__data__0__anchor__in,
	input branch_14__sink_9__data__0__anchor__in,
	input fork_32__branch_13__data__0__anchor__in,
	input branch_18__phi_42__ready__0__anchor__in,
	input fork_34__branch_21__data__0__anchor__in,
	input branch_2__sink_2__valid__0__anchor__in,
	input [31 : 0] branch_36__phi_82__data__0__anchor__in,
	input [31 : 0] Buffer_19__phi_n1__data__0__anchor__in,
	input phi_n12__store_1__ready__0__anchor__in,
	input [31 : 0] phi_n27__fork_28__data__0__anchor__in,
	input Buffer_8__phi_82__ready__0__anchor__in,
	input cst_11__add_54__valid__0__anchor__in,
	input cst_25__MC_A__ready__0__anchor__in,
	input fork_41__branch_42__valid__0__anchor__in,
	input start_0__forkC_44__data__0__anchor__in,
	input mul_89__mul_93__valid__0__anchor__in,
	input [31 : 0] phi_n12__store_1__data__0__anchor__in,
	input phiC_41__ret_0__data__0__anchor__in,
	input branch_6__sink_6__ready__0__anchor__in,
	input phiC_30__branchC_49__data__0__anchor__in,
	input phiC_29__phi_3__valid__0__anchor__in,
	input cst_0__branch_0__ready__0__anchor__in,
	input fork_30__branchC_47__ready__0__anchor__in,
	input forkC_54__brCst_block11__data__0__anchor__in,
	input Buffer_7__phiC_36__valid__0__anchor__in,
	input brCst_block12__fork_40__ready__0__anchor__in,
	input beta__branch_1__valid__0__anchor__in,
	input fork_39__branchC_56__valid__0__anchor__in,
	input branchC_49__Buffer_16__data__0__anchor__in,
	input phiC_39__fork_65__ready__0__anchor__in,
	input fork_11__add_85__valid__0__anchor__in,
	input fork_37__branchC_54__ready__0__anchor__in,
	input phi_77__fork_10__ready__0__anchor__in,
	input branch_34__phi_77__ready__0__anchor__in,
	input phi_n9__branch_16__valid__0__anchor__in,
	input [5 : 0] branch_7__sink_7__data__0__anchor__in,
	input branch_32__sink_22__valid__0__anchor__in,
	input fork_8__store_2__ready__0__anchor__in,
	input [2 : 0] source_13__cst_20__data__0__anchor__in,
	input branch_12__phi_n8__valid__0__anchor__in,
	input branch_0__sink_0__ready__0__anchor__in,
	input forkC_48__branchC_50__valid__0__anchor__in,
	input [5 : 0] add_100__fork_14__data__0__anchor__in,
	input fork_8__load_66__valid__0__anchor__in,
	input forkC_54__cst_18__data__0__anchor__in,
	input [5 : 0] branch_18__phi_42__data__0__anchor__in,
	input forkC_49__cst_9__data__0__anchor__in,
	input phiC_32__phi_36__valid__0__anchor__in,
	input add_94__branch_40__ready__0__anchor__in,
	input forkC_53__cst_27__ready__0__anchor__in,
	input branch_24__phi_n13__ready__0__anchor__in,
	input load_22__MC_v2__valid__0__anchor__in,
	input fork_23__branch_25__ready__0__anchor__in,
	input cst_11__add_54__ready__0__anchor__in,
	input fork_34__branch_19__data__0__anchor__in,
	input branchC_48__Buffer_20__data__0__anchor__in,
	input branch_0__sink_0__valid__0__anchor__in,
	input load_14__MC_v1__valid__0__anchor__in,
	input branch_5__phi_n6__ready__0__anchor__in,
	input branch_18__sink_13__ready__0__anchor__in,
	input load_19__MC_u2__ready__0__anchor__in,
	input [31 : 0] branch_2__sink_2__data__0__anchor__in,
	input [5 : 0] store_2__MC_x__data__1__anchor__in,
	input fork_36__branch_28__ready__0__anchor__in,
	input forkC_46__cst_25__data__0__anchor__in,
	input add_53__branch_22__ready__0__anchor__in,
	input branch_34__sink_23__ready__0__anchor__in,
	input phiC_28__phi_1__ready__0__anchor__in,
	input [31 : 0] phi_n25__branch_44__data__0__anchor__in,
	input [31 : 0] phi_n3__branch_12__data__0__anchor__in,
	input [5 : 0] branch_39__phi_n26__data__0__anchor__in,
	input fork_17__shl_4__valid__0__anchor__in,
	input forkC_46__cst_25__valid__0__anchor__in,
	input branch_17__phi_41__valid__0__anchor__in,
	input forkC_44__brCst_block1__data__0__anchor__in,
	input fork_26__add_100__valid__0__anchor__in,
	input branch_22__phi_n12__valid__0__anchor__in,
	input [31 : 0] branch_40__phi_n23__data__0__anchor__in,
	input forkC_48__cst_8__data__0__anchor__in,
	input fork_31__branch_10__valid__0__anchor__in,
	input fork_1__icmp_30__ready__0__anchor__in,
	input [5 : 0] fork_20__add_59__data__0__anchor__in,
	input branch_30__sink_20__ready__0__anchor__in,
	input Buffer_0__phi_77__ready__0__anchor__in,
	input phi_n18__branch_26__valid__0__anchor__in,
	input forkC_57__cst_28__ready__0__anchor__in,
	input branch_0__sink_0__data__0__anchor__in,
	input branch_44__Buffer_11__valid__0__anchor__in,
	input phiC_35__forkC_52__ready__0__anchor__in,
	input [5 : 0] store_1__MC_x__data__1__anchor__in,
	input forkC_45__cst_1__valid__0__anchor__in,
	input [31 : 0] phi_n23__store_3__data__0__anchor__in,
	input fork_22__add_44__valid__0__anchor__in,
	input fork_41__branchC_58__valid__0__anchor__in,
	input [31 : 0] branch_29__Buffer_24__data__0__anchor__in,
	input fork_29__branch_1__valid__0__anchor__in,
	input [5 : 0] Buffer_15__phi_n26__data__0__anchor__in,
	input [5 : 0] load_14__MC_v1__data__0__anchor__in,
	input fork_40__branch_38__valid__0__anchor__in,
	input phiC_33__fork_62__ready__0__anchor__in,
	input beta__branch_1__ready__0__anchor__in,
	input fork_11__load_92__ready__0__anchor__in,
	input branch_27__sink_18__valid__0__anchor__in,
	input forkC_53__branchC_55__data__0__anchor__in,
	input branchC_54__sink_36__ready__0__anchor__in,
	input MC_u2__end_0__valid__0__anchor__in,
	input phi_n16__fork_22__ready__0__anchor__in,
	input fork_40__branchC_57__ready__0__anchor__in,
	input mul_48__mul_52__valid__0__anchor__in,
	input branch_27__sink_18__ready__0__anchor__in,
	input source_7__cst_11__data__0__anchor__in,
	input branchC_55__phiC_37__ready__0__anchor__in,
	input phi_n27__fork_28__ready__0__anchor__in,
	input fork_34__branchC_51__ready__0__anchor__in,
	input [31 : 0] phi_n20__branch_33__data__0__anchor__in,
	input fork_30__branch_3__ready__0__anchor__in,
	input phi_n22__branch_38__ready__0__anchor__in,
	input forkC_54__cst_18__valid__0__anchor__in,
	input fork_37__branch_31__ready__0__anchor__in,
	input MC_u2__end_0__data__0__anchor__in,
	input source_14__cst_21__valid__0__anchor__in,
	input fork_30__branch_3__valid__0__anchor__in,
	input [31 : 0] fork_23__branch_25__data__0__anchor__in,
	input Buffer_20__phiC_29__ready__0__anchor__in,
	input phi_83__fork_11__valid__0__anchor__in,
	input [5 : 0] branch_7__Buffer_25__data__0__anchor__in,
	input phiC_38__phi_77__valid__0__anchor__in,
	input [31 : 0] MC_A__load_8__data__0__anchor__in,
	input branchC_46__sink_32__ready__0__anchor__in,
	input fork_31__branch_10__data__0__anchor__in,
	input load_11__mul_15__valid__0__anchor__in,
	input load_22__MC_v2__ready__0__anchor__in,
	input fork_41__branch_40__valid__0__anchor__in,
	input forkC_44__branchC_46__data__0__anchor__in,
	input forkC_55__brCst_block12__valid__0__anchor__in,
	input cst_27__MC_x__ready__0__anchor__in,
	input branch_29__phi_n19__valid__0__anchor__in,
	input Buffer_20__phiC_29__data__0__anchor__in,
	input load_69__add_70__ready__0__anchor__in,
	input branchC_58__phiC_40__data__0__anchor__in,
	input branchC_46__phiC_28__valid__0__anchor__in,
	input source_5__cst_7__ready__0__anchor__in,
	input [31 : 0] alpha__branch_2__data__0__anchor__in,
	input forkC_44__branchC_46__valid__0__anchor__in,
	input [31 : 0] Buffer_30__forkC_55__data__0__anchor__in,
	input cst_23__add_100__valid__0__anchor__in,
	input branch_27__Buffer_13__valid__0__anchor__in,
	input forkC_53__branchC_55__valid__0__anchor__in,
	input forkC_48__branchC_50__ready__0__anchor__in,
	input [31 : 0] load_47__mul_48__data__0__anchor__in,
	input [31 : 0] y_din1,
	input [5 : 0] add_73__fork_9__data__0__anchor__in,
	input phiC_30__branchC_49__valid__0__anchor__in,
	input [31 : 0] u2_din1,
	input [5 : 0] phi_3__fork_0__data__0__anchor__in,
	input add_26__store_0__ready__0__anchor__in,
	input load_19__MC_u2__valid__0__anchor__in,
	input branch_6__phi_n7__valid__0__anchor__in,
	input ret_0__end_0__valid__0__anchor__in,
	input branchC_52__Buffer_21__valid__0__anchor__in,
	input [5 : 0] fork_7__icmp_60__data__0__anchor__in,
	input fork_32__branchC_49__ready__0__anchor__in,
	input [31 : 0] MC_v2__load_22__data__0__anchor__in,
	input MC_u1__load_11__ready__0__anchor__in,
	input MC_z__end_0__data__0__anchor__in,
	input [5 : 0] cst_21__add_95__data__0__anchor__in,
	input [5 : 0] fork_1__icmp_30__data__0__anchor__in,
	input cst_14__icmp_60__ready__0__anchor__in,
	input [5 : 0] fork_0__load_14__data__0__anchor__in,
	input cst_1__branch_3__data__0__anchor__in,
	input [5 : 0] branch_42__phi_n24__data__0__anchor__in,
	input start_0__forkC_44__valid__0__anchor__in,
	input [31 : 0] branch_13__phi_n9__data__0__anchor__in,
	input phi_63__fork_8__ready__0__anchor__in,
	input phi_n4__branch_13__valid__0__anchor__in,
	input branch_42__phi_n24__valid__0__anchor__in,
	input fork_20__add_59__ready__0__anchor__in,
	input phiC_30__branchC_49__ready__0__anchor__in,
	input [31 : 0] v1_din1,
	input forkC_51__branchC_53__valid__0__anchor__in,
	input branchC_52__phiC_34__ready__0__anchor__in,
	input cst_8__branch_14__data__0__anchor__in,
	input fork_35__branch_26__ready__0__anchor__in,
	input fork_4__load_51__valid__0__anchor__in,
	input Buffer_27__phiC_32__ready__0__anchor__in,
	input load_69__MC_z__ready__0__anchor__in,
	input MC_w__end_0__data__0__anchor__in,
	input MC_z__end_0__ready__0__anchor__in,
	input [31 : 0] cst_27__MC_x__data__0__anchor__in,
	input branchC_46__phiC_28__data__0__anchor__in,
	input branch_42__phi_n24__ready__0__anchor__in,
	input phiC_34__forkC_51__ready__0__anchor__in,
	input forkC_51__cst_26__data__0__anchor__in,
	input fork_39__branch_34__data__0__anchor__in,
	input cst_28__MC_w__valid__0__anchor__in,
	input phiC_32__phi_36__ready__0__anchor__in,
	input phiC_29__phi_3__ready__0__anchor__in,
	input branch_23__Buffer_3__valid__0__anchor__in,
	input [5 : 0] branch_8__Buffer_14__data__0__anchor__in,
	input cst_19__branch_37__ready__0__anchor__in,
	input forkC_48__cst_8__valid__0__anchor__in,
	input forkC_48__cst_8__ready__0__anchor__in,
	input branch_14__sink_9__valid__0__anchor__in,
	input branchC_50__sink_34__valid__0__anchor__in,
	input [11 : 0] load_8__MC_A__data__0__anchor__in,
	input phiC_29__forkC_46__valid__0__anchor__in,
	input branch_34__phi_77__valid__0__anchor__in,
	input fork_65__phi_83__valid__0__anchor__in,
	input forkC_46__branchC_48__data__0__anchor__in,
	input branchC_51__phiC_33__data__0__anchor__in,
	input fork_37__branchC_54__data__0__anchor__in,
	input MC_v2__end_0__ready__0__anchor__in,
	input branch_41__sink_29__ready__0__anchor__in,
	input branch_29__Buffer_24__ready__0__anchor__in,
	input forkC_49__branchC_51__valid__0__anchor__in,
	input fork_1__branch_7__ready__0__anchor__in,
	input phi_3__fork_0__valid__0__anchor__in,
	input branch_40__Buffer_8__valid__0__anchor__in,
	input fork_38__branch_33__valid__0__anchor__in,
	input fork_39__branch_34__ready__0__anchor__in,
	input [5 : 0] fork_8__store_2__data__0__anchor__in,
	input phiC_28__phi_1__data__0__anchor__in,
	input Buffer_4__phi_n6__valid__0__anchor__in,
	input [31 : 0] cst_25__MC_A__data__0__anchor__in,
	input source_13__cst_20__valid__0__anchor__in,
	input fork_29__branch_2__valid__0__anchor__in,
	input Buffer_23__phi_n27__valid__0__anchor__in,
	input [31 : 0] branch_44__Buffer_11__data__0__anchor__in,
	input Buffer_16__phiC_28__valid__0__anchor__in,
	input phi_n24__fork_26__ready__0__anchor__in,
	input branchC_49__phiC_31__valid__0__anchor__in,
	input fork_34__branchC_51__valid__0__anchor__in,
	input branch_19__phi_n17__ready__0__anchor__in,
	input mul_15__add_16__valid__0__anchor__in,
	input forkC_53__cst_27__valid__0__anchor__in,
	input branch_15__sink_10__ready__0__anchor__in,
	input load_11__mul_15__ready__0__anchor__in,
	input cst_9__branch_18__data__0__anchor__in,
	input fork_34__branch_17__data__0__anchor__in,
	input fork_29__branchC_46__ready__0__anchor__in,
	input cst_3__shl_25__ready__0__anchor__in,
	input load_47__mul_48__valid__0__anchor__in,
	input cst_19__branch_37__valid__0__anchor__in,
	input [5 : 0] fork_10__branch_39__data__0__anchor__in,
	input branchC_55__phiC_37__data__0__anchor__in,
	input icmp_30__fork_31__valid__0__anchor__in,
	input forkC_45__brCst_block2__valid__0__anchor__in,
	input fork_13__branch_41__valid__0__anchor__in,
	input fork_62__phi_42__ready__0__anchor__in,
	input [31 : 0] phi_n22__branch_38__data__0__anchor__in,
	input source_15__cst_22__ready__0__anchor__in,
	input load_80__branch_36__ready__0__anchor__in,
	input branch_32__Buffer_10__ready__0__anchor__in,
	input [31 : 0] branch_25__phi_n14__data__0__anchor__in,
	input fork_32__branch_12__ready__0__anchor__in,
	input MC_x__load_39__ready__0__anchor__in,
	input [5 : 0] Buffer_25__phi_3__data__0__anchor__in,
	input source_1__cst_3__valid__0__anchor__in,
	input phi_n10__branch_19__valid__0__anchor__in,
	input fork_32__branchC_49__data__0__anchor__in,
	input branchC_48__phiC_30__data__0__anchor__in,
	input [11 : 0] fork_11__add_85__data__0__anchor__in,
	input source_10__cst_14__valid__0__anchor__in,
	input fork_29__branch_2__data__0__anchor__in,
	input Buffer_11__phi_n22__valid__0__anchor__in,
	input cst_1__branch_3__ready__0__anchor__in,
	input [31 : 0] branch_33__Buffer_28__data__0__anchor__in,
	input branchC_49__phiC_31__data__0__anchor__in,
	input [31 : 0] w_din1,
	input phi_n26__fork_27__ready__0__anchor__in,
	input phi_n13__fork_20__valid__0__anchor__in,
	input branch_41__sink_29__valid__0__anchor__in,
	input shl_4__add_5__ready__0__anchor__in,
	input fork_34__branchC_51__data__0__anchor__in,
	input MC_w__load_80__valid__0__anchor__in,
	input [31 : 0] branch_22__Buffer_12__data__0__anchor__in,
	input branchC_49__phiC_31__ready__0__anchor__in,
	input Buffer_18__phi_n18__valid__0__anchor__in,
	input add_24__store_0__valid__0__anchor__in,
	input [31 : 0] beta_din,
	input branch_9__Buffer_4__valid__0__anchor__in,
	input MC_y__end_0__ready__0__anchor__in,
	input ret_0__end_0__data__0__anchor__in,
	input branch_19__phi_n17__valid__0__anchor__in,
	input branch_33__Buffer_28__valid__0__anchor__in,
	input MC_y__load_51__valid__0__anchor__in,
	input branch_36__sink_25__ready__0__anchor__in,
	input fork_31__branch_10__ready__0__anchor__in,
	input branch_35__sink_24__ready__0__anchor__in,
	input forkC_52__branchC_54__valid__0__anchor__in,
	input fork_41__branch_42__data__0__anchor__in,
	input MC_u2__end_0__ready__0__anchor__in,
	input add_70__store_2__ready__0__anchor__in,
	input [5 : 0] fork_14__branch_45__data__0__anchor__in,
	input [31 : 0] cst_28__MC_w__data__0__anchor__in,
	input phi_n23__store_3__valid__0__anchor__in,
	input forkC_49__cst_9__valid__0__anchor__in,
	input cst_1__branch_3__valid__0__anchor__in,
	input fork_37__branch_30__data__0__anchor__in,
	input fork_35__branchC_52__valid__0__anchor__in,
	input branch_14__phi_36__valid__0__anchor__in,
	input branch_17__sink_12__valid__0__anchor__in,
	input Buffer_22__phi_n17__ready__0__anchor__in,
	input fork_14__icmp_101__ready__0__anchor__in,
	input branch_25__phi_n14__ready__0__anchor__in,
	input branch_44__Buffer_11__ready__0__anchor__in,
	input branch_37__phi_83__ready__0__anchor__in,
	input branch_45__Buffer_0__ready__0__anchor__in,
	input phi_n25__branch_44__valid__0__anchor__in,
	input forkC_54__brCst_block11__ready__0__anchor__in,
	input cst_5__icmp_30__ready__0__anchor__in,
	input [5 : 0] branch_39__sink_28__data__0__anchor__in,
	input phi_83__fork_11__ready__0__anchor__in,
	input forkC_45__brCst_block2__ready__0__anchor__in,
	input phiC_29__phi_3__data__0__anchor__in,
	input branch_41__Buffer_29__ready__0__anchor__in,
	input fork_41__branch_43__ready__0__anchor__in,
	input cst_21__add_95__valid__0__anchor__in,
	input branch_24__phi_n13__valid__0__anchor__in,
	input branchC_53__Buffer_27__valid__0__anchor__in,
	input fork_17__load_11__valid__0__anchor__in,
	input add_100__fork_14__ready__0__anchor__in,
	input [5 : 0] add_54__fork_6__data__0__anchor__in,
	input brCst_block11__fork_39__valid__0__anchor__in,
	input fork_35__branch_22__data__0__anchor__in,
	input fork_65__phi_83__data__0__anchor__in,
	input [31 : 0] branch_2__phi_n1__data__0__anchor__in,
	input fork_30__branch_4__valid__0__anchor__in,
	input branchC_55__phiC_37__valid__0__anchor__in,
	input phiC_37__forkC_54__ready__0__anchor__in,
	input [31 : 0] phi_n21__branch_35__data__0__anchor__in,
	input icmp_101__fork_42__valid__0__anchor__in,
	input [5 : 0] phi_n16__fork_22__data__0__anchor__in,
	input fork_22__add_44__ready__0__anchor__in,
	input fork_42__branchC_59__data__0__anchor__in,
	input branchC_54__phiC_36__data__0__anchor__in,
	input load_51__MC_y__ready__0__anchor__in,
	input fork_65__phi_82__valid__0__anchor__in,
	input [5 : 0] source_3__cst_5__data__0__anchor__in,
	input phiC_39__branchC_58__data__0__anchor__in,
	input Buffer_13__phi_n10__valid__0__anchor__in,
	input Buffer_0__phi_77__valid__0__anchor__in,
	input Buffer_21__phiC_33__ready__0__anchor__in,
	input [5 : 0] fork_17__load_19__data__0__anchor__in,
	input branch_20__sink_15__valid__0__anchor__in,
	input branchC_51__phiC_33__ready__0__anchor__in,
	input branchC_57__sink_38__valid__0__anchor__in,
	input end_ready,
	input fork_32__branch_11__valid__0__anchor__in,
	input phi_n14__branch_27__ready__0__anchor__in,
	input [31 : 0] phi_41__add_53__data__0__anchor__in,
	input Buffer_30__forkC_55__valid__0__anchor__in,
	input branchC_51__phiC_33__valid__0__anchor__in,
	input branch_2__phi_n1__valid__0__anchor__in,
	input branch_11__sink_8__ready__0__anchor__in,
	input branch_36__phi_82__ready__0__anchor__in,
	input forkC_51__cst_26__ready__0__anchor__in,
	input phiC_39__fork_65__data__0__anchor__in,
	input [31 : 0] MC_w__load_80__data__0__anchor__in,
	input fork_33__branchC_50__data__0__anchor__in,
	input [31 : 0] branch_9__phi_n3__data__0__anchor__in,
	input fork_28__mul_89__ready__0__anchor__in,
	input fork_4__shl_43__ready__0__anchor__in,
	input fork_42__branch_44__ready__0__anchor__in,
	input branch_39__phi_n26__valid__0__anchor__in,
	input [5 : 0] branch_23__sink_17__data__0__anchor__in,
	input fork_0__add_26__ready__0__anchor__in,
	input icmp_55__fork_35__data__0__anchor__in,
	input phi_n10__branch_19__ready__0__anchor__in,
	input branch_16__phi_n11__valid__0__anchor__in,
	input [31 : 0] MC_v1__load_14__data__0__anchor__in,
	input branchC_56__phiC_38__data__0__anchor__in,
	input fork_14__branch_45__ready__0__anchor__in,
	input fork_20__store_1__ready__0__anchor__in,
	input alpha__branch_2__valid__0__anchor__in,
	input forkC_48__brCst_block5__data__0__anchor__in,
	input phi_63__fork_8__valid__0__anchor__in,
	input [31 : 0] x_din0,
	input fork_39__branch_35__valid__0__anchor__in,
	input MC_A__load_88__valid__0__anchor__in,
	input [10 : 0] fork_17__shl_25__data__0__anchor__in,
	input [31 : 0] load_11__mul_15__data__0__anchor__in,
	input [5 : 0] source_5__cst_7__data__0__anchor__in,
	input [31 : 0] load_19__mul_23__data__0__anchor__in,
	input store_1__MC_x__ready__1__anchor__in,
	input branchC_56__phiC_38__valid__0__anchor__in,
	input [31 : 0] add_16__add_24__data__0__anchor__in,
	input fork_33__branch_14__ready__0__anchor__in,
	input [31 : 0] branch_25__Buffer_22__data__0__anchor__in,
	input phi_77__fork_10__valid__0__anchor__in,
	input fork_8__load_69__ready__0__anchor__in,
	input [31 : 0] mul_15__add_16__data__0__anchor__in,
	input branchC_57__phiC_39__ready__0__anchor__in,
	input branch_2__sink_2__ready__0__anchor__in,
	input source_3__cst_5__ready__0__anchor__in,
	input fork_2__icmp_33__valid__0__anchor__in,
	input branch_43__phi_n25__ready__0__anchor__in,
	input source_11__cst_16__ready__0__anchor__in,
	input load_14__mul_15__valid__0__anchor__in,
	input load_14__MC_v1__ready__0__anchor__in,
	input fork_34__branch_21__valid__0__anchor__in,
	input fork_2__icmp_33__ready__0__anchor__in,
	input fork_41__branch_41__data__0__anchor__in,
	input fork_42__branchC_59__ready__0__anchor__in,
	input fork_9__icmp_74__valid__0__anchor__in,
	input phiC_38__Buffer_30__valid__0__anchor__in,
	input [5 : 0] phi_77__fork_10__data__0__anchor__in,
	input [31 : 0] phi_n4__branch_13__data__0__anchor__in,
	input fork_0__load_22__valid__0__anchor__in,
	input [11 : 0] add_85__load_88__data__0__anchor__in,
	input fork_33__branch_14__data__0__anchor__in,
	input [31 : 0] branch_43__phi_n25__data__0__anchor__in,
	input Buffer_29__phi_83__ready__0__anchor__in,
	input fork_33__branch_16__valid__0__anchor__in,
	input add_73__fork_9__ready__0__anchor__in,
	input branchC_47__sink_33__ready__0__anchor__in,
	input [5 : 0] Buffer_3__phi_42__data__0__anchor__in,
	input [5 : 0] branch_30__phi_63__data__0__anchor__in,
	input [5 : 0] branch_24__Buffer_17__data__0__anchor__in,
	input [31 : 0] load_66__add_70__data__0__anchor__in,
	input MC_v2__end_0__valid__0__anchor__in,
	input cst_13__add_59__ready__0__anchor__in,
	input [5 : 0] fork_8__load_69__data__0__anchor__in,
	input [5 : 0] branch_23__Buffer_3__data__0__anchor__in,
	input fork_9__icmp_74__ready__0__anchor__in,
	input branchC_50__phiC_32__data__0__anchor__in,
	input branch_45__sink_31__valid__0__anchor__in,
	input phi_n2__add_32__valid__0__anchor__in,
	input branch_20__phi_n18__valid__0__anchor__in,
	input alpha__branch_2__ready__0__anchor__in,
	input source_17__cst_24__ready__0__anchor__in,
	input forkC_52__cst_15__valid__0__anchor__in,
	input phi_n1__branch_6__ready__0__anchor__in,
	input phi_82__add_94__valid__0__anchor__in,
	input [31 : 0] phi_n11__branch_20__data__0__anchor__in,
	input branch_30__sink_20__valid__0__anchor__in,
	input load_47__MC_A__valid__0__anchor__in,
	input branch_34__sink_23__valid__0__anchor__in,
	input fork_30__branch_5__valid__0__anchor__in,
	input phi_n12__store_1__valid__0__anchor__in,
	input MC_v1__end_0__valid__0__anchor__in,
	input phi_n15__branch_29__valid__0__anchor__in,
	input fork_33__branch_15__data__0__anchor__in,
	input [5 : 0] fork_26__add_100__data__0__anchor__in,
	input fork_8__load_66__ready__0__anchor__in,
	input Buffer_20__phiC_29__valid__0__anchor__in,
	input [5 : 0] fork_17__branch_8__data__0__anchor__in,
	input source_7__cst_11__valid__0__anchor__in,
	input branchC_52__Buffer_21__data__0__anchor__in,
	input MC_v1__load_14__valid__0__anchor__in,
	input load_66__add_70__ready__0__anchor__in,
	input [31 : 0] branch_13__Buffer_19__data__0__anchor__in,
	input fork_17__shl_4__ready__0__anchor__in,
	input fork_17__load_19__ready__0__anchor__in,
	input fork_28__mul_89__valid__0__anchor__in,
	input MC_v1__end_0__data__0__anchor__in,
	input [31 : 0] phi_n0__branch_5__data__0__anchor__in,
	input fork_39__branch_34__valid__0__anchor__in,
	input branchC_55__Buffer_7__valid__0__anchor__in,
	input [31 : 0] branch_16__phi_n11__data__0__anchor__in,
	input store_1__MC_x__valid__0__anchor__in,
	input forkC_54__cst_18__ready__0__anchor__in,
	input Buffer_28__phi_n20__valid__0__anchor__in,
	input source_2__cst_4__ready__0__anchor__in,
	input fork_42__branch_45__ready__0__anchor__in,
	input cst_6__add_32__valid__0__anchor__in,
	input fork_30__branch_5__data__0__anchor__in,
	input Buffer_21__phiC_33__valid__0__anchor__in,
	input store_2__MC_x__ready__1__anchor__in,
	input cst_12__icmp_55__valid__0__anchor__in,
	input fork_40__branch_39__valid__0__anchor__in,
	input forkC_44__cst_0__data__0__anchor__in,
	input [10 : 0] fork_4__shl_43__data__0__anchor__in,
	input [31 : 0] branch_40__Buffer_8__data__0__anchor__in,
	input [31 : 0] add_53__branch_22__data__0__anchor__in,
	input MC_A__end_0__data__0__anchor__in,
	input branchC_48__Buffer_20__ready__0__anchor__in,
	input forkC_46__cst_25__ready__0__anchor__in,
	input fork_35__branch_22__valid__0__anchor__in,
	input [31 : 0] MC_u1__load_11__data__0__anchor__in,
	input brCst_block6__fork_34__data__0__anchor__in,
	input [31 : 0] MC_y__load_51__data__0__anchor__in,
	input MC_A__load_47__valid__0__anchor__in,
	input mul_93__add_94__ready__0__anchor__in,
	input brCst_block12__fork_40__data__0__anchor__in,
	input [5 : 0] fork_27__branch_42__data__0__anchor__in,
	input [5 : 0] branch_42__Buffer_15__data__0__anchor__in,
	input phi_n13__fork_20__ready__0__anchor__in,
	input branch_36__sink_25__valid__0__anchor__in,
	input MC_w__end_0__valid__0__anchor__in,
	input phiC_41__ret_0__ready__0__anchor__in,
	input [5 : 0] add_29__fork_1__data__0__anchor__in,
	input branchC_54__sink_36__valid__0__anchor__in,
	input [5 : 0] fork_4__add_54__data__0__anchor__in,
	input phi_n7__branch_10__valid__0__anchor__in,
	input phiC_33__branchC_52__data__0__anchor__in,
	input fork_36__branchC_53__data__0__anchor__in,
	input fork_42__branch_44__valid__0__anchor__in,
	input phi_n21__branch_35__ready__0__anchor__in,
	input fork_10__load_80__ready__0__anchor__in,
	input phi_42__fork_4__ready__0__anchor__in,
	input load_66__MC_x__ready__0__anchor__in,
	input [5 : 0] branch_37__phi_83__data__0__anchor__in,
	input fork_27__shl_84__valid__0__anchor__in,
	input cst_26__MC_x__ready__0__anchor__in,
	input Buffer_3__phi_42__ready__0__anchor__in,
	input branchC_47__sink_33__valid__0__anchor__in,
	input fork_30__branch_4__ready__0__anchor__in,
	input add_70__store_2__valid__0__anchor__in,
	input fork_41__branchC_58__ready__0__anchor__in,
	input branch_21__phi_n16__ready__0__anchor__in,
	input fork_35__branch_23__data__0__anchor__in,
	input branch_8__Buffer_14__ready__0__anchor__in,
	input add_95__fork_13__valid__0__anchor__in,
	input load_92__mul_93__ready__0__anchor__in,
	input MC_A__load_47__ready__0__anchor__in,
	input fork_62__phi_41__valid__0__anchor__in,
	input [5 : 0] add_59__fork_7__data__0__anchor__in,
	input fork_33__branch_14__valid__0__anchor__in,
	input MC_x__load_92__valid__0__anchor__in,
	input [10 : 0] fork_27__shl_84__data__0__anchor__in,
	input [5 : 0] Buffer_9__phi_36__data__0__anchor__in,
	input Buffer_19__phi_n1__valid__0__anchor__in,
	input forkC_44__brCst_block1__valid__0__anchor__in,
	input phiC_33__fork_62__data__0__anchor__in,
	input phi_n24__fork_26__valid__0__anchor__in,
	input [5 : 0] phi_n2__add_32__data__0__anchor__in,
	input branch_27__Buffer_13__ready__0__anchor__in,
	input [31 : 0] Buffer_12__phi_41__data__0__anchor__in,
	input branch_20__phi_n18__ready__0__anchor__in,
	input Buffer_2__phiC_39__valid__0__anchor__in,
	input [31 : 0] store_0__MC_A__data__0__anchor__in,
	input fork_2__branch_11__valid__0__anchor__in,
	input [5 : 0] cst_17__icmp_74__data__0__anchor__in,
	input brCst_block1__fork_29__valid__0__anchor__in,
	input icmp_74__fork_38__valid__0__anchor__in,
	input branch_8__phi_n2__valid__0__anchor__in,
	input fork_34__branch_18__data__0__anchor__in,
	input source_16__cst_23__data__0__anchor__in,
	input add_85__load_88__ready__0__anchor__in,
	input [5 : 0] phi_n5__fork_17__data__0__anchor__in,
	input fork_35__branch_26__data__0__anchor__in,
	input brCst_block11__fork_39__ready__0__anchor__in,
	input [31 : 0] branch_35__sink_24__data__0__anchor__in,
	input phiC_35__forkC_52__data__0__anchor__in,
	input fork_22__branch_24__ready__0__anchor__in,
	input fork_41__branch_41__ready__0__anchor__in,
	input [31 : 0] add_70__store_2__data__0__anchor__in,
	input phiC_33__fork_62__valid__0__anchor__in,
	input fork_6__branch_23__ready__0__anchor__in,
	input branch_22__Buffer_12__valid__0__anchor__in,
	input Buffer_1__phi_n0__valid__0__anchor__in,
	input phiC_33__branchC_52__valid__0__anchor__in,
	input branchC_52__Buffer_21__ready__0__anchor__in,
	input fork_62__phi_42__data__0__anchor__in,
	input forkC_44__cst_0__valid__0__anchor__in,
	input fork_37__branchC_54__valid__0__anchor__in,
	input branch_28__Buffer_9__ready__0__anchor__in,
	input mul_52__add_53__ready__0__anchor__in,
	input forkC_55__brCst_block12__data__0__anchor__in,
	input MC_A__end_0__valid__0__anchor__in,
	input [5 : 0] add_95__fork_13__data__0__anchor__in,
	input [31 : 0] branch_26__phi_n15__data__0__anchor__in,
	input load_88__MC_A__ready__0__anchor__in,
	input fork_31__branch_8__ready__0__anchor__in,
	input branchC_50__sink_34__data__0__anchor__in,
	input source_0__cst_2__valid__0__anchor__in,
	input fork_27__branch_42__valid__0__anchor__in,
	input [11 : 0] shl_25__add_26__data__0__anchor__in,
	input fork_39__branch_35__ready__0__anchor__in,
	input icmp_101__fork_42__data__0__anchor__in,
	input fork_41__branch_40__ready__0__anchor__in,
	input [31 : 0] v2_din0,
	input fork_8__add_73__valid__0__anchor__in,
	input load_66__add_70__valid__0__anchor__in,
	input brCst_block11__fork_39__data__0__anchor__in,
	input fork_29__branch_0__data__0__anchor__in,
	input cst_22__icmp_96__valid__0__anchor__in,
	input fork_31__branchC_48__valid__0__anchor__in,
	input fork_4__load_51__ready__0__anchor__in,
	input source_10__cst_14__ready__0__anchor__in,
	input icmp_30__fork_31__data__0__anchor__in,
	input load_11__MC_u1__ready__0__anchor__in,
	input [31 : 0] fork_28__mul_89__data__0__anchor__in,
	input fork_36__branch_29__valid__0__anchor__in,
	input load_51__mul_52__valid__0__anchor__in,
	input [5 : 0] fork_3__load_39__data__0__anchor__in,
	input [5 : 0] cst_4__add_29__data__0__anchor__in,
	input branchC_58__Buffer_2__valid__0__anchor__in,
	input forkC_52__branchC_54__data__0__anchor__in,
	input Buffer_27__phiC_32__data__0__anchor__in,
	input branch_32__sink_22__ready__0__anchor__in,
	input [31 : 0] phi_82__add_94__data__0__anchor__in,
	input [5 : 0] fork_9__icmp_74__data__0__anchor__in,
	input brCst_block12__fork_40__valid__0__anchor__in,
	input [31 : 0] Buffer_22__phi_n17__data__0__anchor__in,
	input branch_14__phi_36__ready__0__anchor__in,
	input [31 : 0] branch_17__sink_12__data__0__anchor__in,
	input fork_40__branch_38__ready__0__anchor__in,
	input cst_6__add_32__ready__0__anchor__in,
	input fork_31__branchC_48__ready__0__anchor__in,
	input branch_22__Buffer_12__ready__0__anchor__in,
	input [31 : 0] load_14__mul_15__data__0__anchor__in,
	input icmp_33__fork_32__ready__0__anchor__in,
	input forkC_48__brCst_block5__ready__0__anchor__in,
	input phi_n3__branch_12__ready__0__anchor__in,
	input phi_n8__branch_15__ready__0__anchor__in,
	input branchC_57__phiC_39__data__0__anchor__in,
	input fork_35__branch_23__ready__0__anchor__in,
	input add_24__store_0__ready__0__anchor__in,
	input source_2__cst_4__data__0__anchor__in,
	input fork_30__branch_4__data__0__anchor__in,
	input [5 : 0] store_3__MC_w__data__1__anchor__in,
	input branchC_56__phiC_38__ready__0__anchor__in,
	input [11 : 0] add_44__load_47__data__0__anchor__in,
	input branch_22__phi_n12__ready__0__anchor__in,
	input cst_8__branch_14__valid__0__anchor__in,
	input branch_25__Buffer_22__valid__0__anchor__in,
	input forkC_49__branchC_51__data__0__anchor__in,
	input icmp_96__fork_41__ready__0__anchor__in,
	input fork_34__branch_20__data__0__anchor__in,
	input [5 : 0] phi_1__branch_4__data__0__anchor__in,
	input fork_29__branch_1__data__0__anchor__in,
	input fork_40__branch_36__data__0__anchor__in,
	input fork_41__branchC_58__data__0__anchor__in,
	input brCst_block1__fork_29__ready__0__anchor__in,
	input brCst_block9__fork_37__ready__0__anchor__in,
	input [5 : 0] cst_7__icmp_33__data__0__anchor__in,
	input fork_36__branch_28__valid__0__anchor__in,
	input [31 : 0] add_94__branch_40__data__0__anchor__in,
	input fork_33__branch_16__data__0__anchor__in,
	input forkC_49__brCst_block6__data__0__anchor__in,
	input source_1__cst_3__ready__0__anchor__in,
	input phi_n1__branch_6__valid__0__anchor__in,
	input [5 : 0] phi_63__fork_8__data__0__anchor__in,
	input branchC_51__sink_35__ready__0__anchor__in,
	input [5 : 0] cst_13__add_59__data__0__anchor__in,
	input fork_3__branch_21__valid__0__anchor__in,
	input MC_z__end_0__valid__0__anchor__in,
	input [31 : 0] branch_38__phi_n27__data__0__anchor__in,
	input branch_30__sink_20__data__0__anchor__in,
	input brCst_block2__fork_30__valid__0__anchor__in,
	input source_9__cst_13__valid__0__anchor__in,
	input MC_x__end_0__data__0__anchor__in,
	input phiC_29__forkC_46__ready__0__anchor__in,
	input branch_1__phi_n0__ready__0__anchor__in,
	input fork_31__branch_7__valid__0__anchor__in,
	input fork_17__branch_8__ready__0__anchor__in,
	input load_8__MC_A__ready__0__anchor__in,
	input fork_65__phi_82__ready__0__anchor__in,
	input fork_6__branch_23__valid__0__anchor__in,
	input [10 : 0] cst_20__shl_84__data__0__anchor__in,
	input fork_13__branch_41__ready__0__anchor__in,
	input fork_14__icmp_101__valid__0__anchor__in,
	input forkC_52__cst_15__data__0__anchor__in,
	input Buffer_2__phiC_39__data__0__anchor__in,
	input brCst_block9__fork_37__valid__0__anchor__in,
	input [5 : 0] fork_6__branch_23__data__0__anchor__in,
	input fork_36__branch_27__data__0__anchor__in,
	input fork_33__branch_15__ready__0__anchor__in,
	input branchC_49__Buffer_16__valid__0__anchor__in,
	input branch_41__Buffer_29__valid__0__anchor__in,
	input [31 : 0] A_din1,
	input brCst_block9__fork_37__data__0__anchor__in,
	input fork_8__load_69__valid__0__anchor__in,
	input forkC_46__branchC_48__valid__0__anchor__in,
	input forkC_46__branchC_48__ready__0__anchor__in,
	input Buffer_19__phi_n1__ready__0__anchor__in,
	input branch_26__phi_n15__ready__0__anchor__in,
	input phi_1__branch_4__ready__0__anchor__in,
	input cst_8__branch_14__ready__0__anchor__in,
	input forkC_54__branchC_56__data__0__anchor__in,
	input phiC_28__forkC_45__data__0__anchor__in,
	input branch_10__phi_n4__valid__0__anchor__in,
	input phi_n5__fork_17__valid__0__anchor__in,
	input add_44__load_47__ready__0__anchor__in,
	input Buffer_5__phi_n7__ready__0__anchor__in,
	input mul_23__add_24__ready__0__anchor__in,
	input source_11__cst_16__valid__0__anchor__in,
	input branch_43__Buffer_23__valid__0__anchor__in,
	input load_8__add_16__ready__0__anchor__in,
	input branch_39__sink_28__ready__0__anchor__in,
	input phiC_41__ret_0__valid__0__anchor__in,
	input phi_42__fork_4__valid__0__anchor__in,
	input Buffer_22__phi_n17__valid__0__anchor__in,
	input phiC_28__forkC_45__valid__0__anchor__in,
	input phiC_40__forkC_57__ready__0__anchor__in,
	input branchC_57__sink_38__ready__0__anchor__in,
	input [31 : 0] phiC_38__Buffer_30__data__0__anchor__in,
	input [31 : 0] Buffer_13__phi_n10__data__0__anchor__in,
	input branchC_54__phiC_36__ready__0__anchor__in,
	input branchC_54__phiC_36__valid__0__anchor__in,
	input phi_n18__branch_26__ready__0__anchor__in,
	input [5 : 0] source_8__cst_12__data__0__anchor__in,
	input Buffer_25__phi_3__ready__0__anchor__in,
	input branchC_48__phiC_30__ready__0__anchor__in,
	input add_95__fork_13__ready__0__anchor__in,
	input [31 : 0] branch_22__phi_n12__data__0__anchor__in,
	input branch_7__sink_7__valid__0__anchor__in,
	input source_12__cst_17__ready__0__anchor__in,
	input phi_41__add_53__valid__0__anchor__in,
	input fork_4__add_54__ready__0__anchor__in,
	input branch_24__Buffer_17__ready__0__anchor__in,
	input forkC_57__branchC_59__data__0__anchor__in,
	input fork_8__store_2__valid__0__anchor__in,
	input MC_x__end_0__ready__0__anchor__in,
	input branch_5__sink_5__ready__0__anchor__in,
	input MC_u1__end_0__data__0__anchor__in,
	input fork_30__branch_6__data__0__anchor__in,
	input branchC_46__sink_32__valid__0__anchor__in,
	input [10 : 0] cst_3__shl_25__data__0__anchor__in,
	input Buffer_21__phiC_33__data__0__anchor__in,
	input branch_38__phi_n27__valid__0__anchor__in,
	input Buffer_15__phi_n26__valid__0__anchor__in,
	input MC_x__load_39__valid__0__anchor__in,
	input [2 : 0] source_0__cst_2__data__0__anchor__in,
	input [5 : 0] branch_11__Buffer_26__data__0__anchor__in,
	input branch_16__sink_11__valid__0__anchor__in,
	input phi_36__fork_3__valid__0__anchor__in,
	input cst_28__MC_w__ready__0__anchor__in,
	input [31 : 0] mul_52__add_53__data__0__anchor__in,
	input branch_4__sink_4__ready__0__anchor__in,
	input phiC_38__Buffer_30__ready__0__anchor__in,
	input phi_n15__branch_29__ready__0__anchor__in,
	input branch_31__sink_21__ready__0__anchor__in,
	input icmp_96__fork_41__data__0__anchor__in,
	input branchC_56__sink_37__ready__0__anchor__in,
	input [5 : 0] cst_24__icmp_101__data__0__anchor__in,
	input mul_23__add_24__valid__0__anchor__in,
	input [5 : 0] branch_14__phi_36__data__0__anchor__in,
	input fork_42__branch_45__valid__0__anchor__in,
	input fork_35__branch_26__valid__0__anchor__in,
	input branch_1__phi_n0__valid__0__anchor__in,
	input branch_33__phi_n21__ready__0__anchor__in,
	input source_16__cst_23__ready__0__anchor__in,
	input fork_29__branchC_46__data__0__anchor__in,
	input store_0__MC_A__valid__1__anchor__in,
	input phiC_31__forkC_48__valid__0__anchor__in,
	input MC_v2__end_0__data__0__anchor__in,
	input fork_35__branch_24__valid__0__anchor__in,
	input store_0__MC_A__ready__0__anchor__in,
	input cst_7__icmp_33__ready__0__anchor__in,
	input add_100__fork_14__valid__0__anchor__in,
	input [5 : 0] branch_11__sink_8__data__0__anchor__in,
	input [31 : 0] branch_20__sink_15__data__0__anchor__in,
	input cst_7__icmp_33__valid__0__anchor__in,
	input forkC_53__cst_27__data__0__anchor__in,
	input MC_u1__end_0__ready__0__anchor__in,
	input [11 : 0] fork_0__add_26__data__0__anchor__in,
	input forkC_55__branchC_57__valid__0__anchor__in,
	input branch_4__phi_n5__valid__0__anchor__in,
	input forkC_45__brCst_block2__data__0__anchor__in,
	input fork_3__load_39__ready__0__anchor__in,
	input [5 : 0] fork_3__branch_21__data__0__anchor__in,
	input cst_10__shl_43__ready__0__anchor__in,
	input [5 : 0] Buffer_0__phi_77__data__0__anchor__in,
	input store_3__MC_w__valid__1__anchor__in,
	input fork_40__branch_36__valid__0__anchor__in,
	input phi_n9__branch_16__ready__0__anchor__in,
	input phiC_38__phi_77__data__0__anchor__in,
	input [11 : 0] shl_43__add_44__data__0__anchor__in,
	input fork_35__branch_25__valid__0__anchor__in,
	input phiC_37__forkC_54__data__0__anchor__in,
	input branch_8__Buffer_14__valid__0__anchor__in,
	input Buffer_11__phi_n22__ready__0__anchor__in,
	input Buffer_5__phi_n7__valid__0__anchor__in,
	input shl_25__add_26__ready__0__anchor__in,
	input branch_39__phi_n26__ready__0__anchor__in,
	input phiC_39__branchC_58__valid__0__anchor__in,
	input phiC_36__forkC_53__valid__0__anchor__in,
	input fork_31__branch_8__valid__0__anchor__in,
	input [5 : 0] branch_28__sink_19__data__0__anchor__in,
	input branch_33__Buffer_28__ready__0__anchor__in,
	input MC_y__load_51__ready__0__anchor__in,
	input [31 : 0] branch_19__phi_n17__data__0__anchor__in,
	input branch_8__phi_n2__ready__0__anchor__in,
	input branchC_51__sink_35__valid__0__anchor__in,
	input branch_20__sink_15__ready__0__anchor__in,
	input cst_27__MC_x__valid__0__anchor__in,
	input fork_33__branchC_50__valid__0__anchor__in,
	input icmp_55__fork_35__ready__0__anchor__in,
	input branchC_50__phiC_32__valid__0__anchor__in,
	input source_7__cst_11__ready__0__anchor__in,
	input icmp_74__fork_38__ready__0__anchor__in,
	input phi_n26__fork_27__valid__0__anchor__in,
	input phiC_28__phi_1__valid__0__anchor__in,
	input [5 : 0] Buffer_26__phi_1__data__0__anchor__in,
	input fork_17__load_19__valid__0__anchor__in,
	input fork_39__branchC_56__ready__0__anchor__in,
	input [31 : 0] alpha_din,
	input phi_n20__branch_33__valid__0__anchor__in,
	input cst_26__MC_x__valid__0__anchor__in,
	input load_88__mul_89__ready__0__anchor__in,
	input fork_40__branch_37__valid__0__anchor__in,
	input [5 : 0] load_80__MC_w__data__0__anchor__in,
	input icmp_30__fork_31__ready__0__anchor__in,
	input phi_n7__branch_10__ready__0__anchor__in,
	input branch_19__sink_14__valid__0__anchor__in,
	input branch_4__phi_n5__ready__0__anchor__in,
	input cst_5__icmp_30__valid__0__anchor__in,
	input phiC_31__forkC_48__data__0__anchor__in,
	input source_5__cst_7__valid__0__anchor__in,
	input fork_32__branch_12__valid__0__anchor__in,
	input branchC_57__sink_38__data__0__anchor__in,
	input [5 : 0] load_19__MC_u2__data__0__anchor__in,
	input cst_17__icmp_74__valid__0__anchor__in,
	input Buffer_17__phi_n16__ready__0__anchor__in,
	input cst_15__branch_30__valid__0__anchor__in,
	input icmp_33__fork_32__data__0__anchor__in,
	input forkC_55__cst_19__data__0__anchor__in,
	input fork_7__icmp_60__valid__0__anchor__in,
	input load_92__MC_x__valid__0__anchor__in,
	input forkC_49__branchC_51__ready__0__anchor__in,
	input fork_9__branch_32__ready__0__anchor__in,
	input branch_45__sink_31__ready__0__anchor__in,
	input branch_45__Buffer_0__valid__0__anchor__in,
	input phiC_32__phi_36__data__0__anchor__in,
	input source_13__cst_20__ready__0__anchor__in,
	input branch_11__sink_8__valid__0__anchor__in,
	input fork_0__add_5__ready__0__anchor__in,
	input branch_35__phi_n22__valid__0__anchor__in,
	input [31 : 0] Buffer_28__phi_n20__data__0__anchor__in,
	input add_32__fork_2__valid__0__anchor__in,
	input branch_12__Buffer_1__valid__0__anchor__in,
	input fork_20__store_1__valid__0__anchor__in,
	input fork_9__branch_32__valid__0__anchor__in,
	input fork_2__branch_11__ready__0__anchor__in,
	input source_9__cst_13__ready__0__anchor__in,
	input [31 : 0] mul_23__add_24__data__0__anchor__in,
	input [5 : 0] cst_5__icmp_30__data__0__anchor__in,
	input phi_n21__branch_35__valid__0__anchor__in,
	input branchC_51__sink_35__data__0__anchor__in,
	input load_39__branch_17__valid__0__anchor__in,
	input [11 : 0] store_0__MC_A__data__1__anchor__in,
	input forkC_57__cst_28__valid__0__anchor__in,
	input mul_93__add_94__valid__0__anchor__in,
	input [5 : 0] load_51__MC_y__data__0__anchor__in,
	input Buffer_10__phi_63__ready__0__anchor__in,
	input phi_n17__fork_23__ready__0__anchor__in,
	input source_9__cst_13__data__0__anchor__in,
	input branch_35__sink_24__valid__0__anchor__in,
	input branch_36__phi_82__valid__0__anchor__in,
	input fork_34__branch_18__valid__0__anchor__in,
	input [5 : 0] cst_12__icmp_55__data__0__anchor__in,
	input source_4__cst_6__valid__0__anchor__in,
	input branchC_48__Buffer_20__valid__0__anchor__in,
	input load_47__mul_48__ready__0__anchor__in,
	input phiC_33__branchC_52__ready__0__anchor__in,
	input [5 : 0] fork_7__branch_28__data__0__anchor__in,
	input [11 : 0] shl_84__add_85__data__0__anchor__in,
	input MC_v2__load_22__ready__0__anchor__in,
	input [5 : 0] fork_26__store_3__data__0__anchor__in,
	input [31 : 0] branch_15__phi_n10__data__0__anchor__in,
	input ret_0__end_0__ready__0__anchor__in,
	input fork_17__shl_25__valid__0__anchor__in,
	input branch_11__Buffer_26__valid__0__anchor__in,
	input icmp_96__fork_41__valid__0__anchor__in,
	input fork_13__icmp_96__valid__0__anchor__in,
	input [5 : 0] fork_8__load_66__data__0__anchor__in,
	input add_32__fork_2__ready__0__anchor__in,
	input fork_38__branch_33__ready__0__anchor__in,
	input [10 : 0] cst_2__shl_4__data__0__anchor__in,
	input [31 : 0] A_din0,
	input Buffer_26__phi_1__ready__0__anchor__in,
	input load_80__MC_w__valid__0__anchor__in,
	input fork_26__add_100__ready__0__anchor__in,
	input [31 : 0] u2_din0,
	input load_14__mul_15__ready__0__anchor__in,
	input fork_1__icmp_30__valid__0__anchor__in,
	input [5 : 0] phi_n26__fork_27__data__0__anchor__in,
	input branchC_58__Buffer_2__ready__0__anchor__in,
	input [31 : 0] MC_x__load_66__data__0__anchor__in,
	input [5 : 0] branch_21__phi_n16__data__0__anchor__in,
	input [31 : 0] branch_10__Buffer_5__data__0__anchor__in,
	input branch_38__sink_27__ready__0__anchor__in,
	input mul_89__mul_93__ready__0__anchor__in,
	input phi_n16__fork_22__valid__0__anchor__in,
	input cst_18__branch_34__valid__0__anchor__in,
	input fork_7__branch_28__valid__0__anchor__in,
	input [5 : 0] branch_24__phi_n13__data__0__anchor__in,
	input add_26__store_0__valid__0__anchor__in,
	input fork_0__load_14__ready__0__anchor__in,
	input [31 : 0] load_8__add_16__data__0__anchor__in,
	input [5 : 0] branch_4__sink_4__data__0__anchor__in,
	input [5 : 0] fork_6__icmp_55__data__0__anchor__in,
	input fork_34__branch_20__ready__0__anchor__in,
	input Buffer_12__phi_41__ready__0__anchor__in,
	input Buffer_14__phi_n5__valid__0__anchor__in,
	input Buffer_16__phiC_28__data__0__anchor__in,
	input load_19__mul_23__ready__0__anchor__in,
	input Buffer_29__phi_83__valid__0__anchor__in,
	input shl_4__add_5__valid__0__anchor__in,
	input [5 : 0] phi_42__fork_4__data__0__anchor__in,
	input branchC_58__Buffer_2__data__0__anchor__in,
	input [11 : 0] shl_4__add_5__data__0__anchor__in,
	input phiC_39__branchC_58__ready__0__anchor__in,
	input [31 : 0] branch_6__phi_n7__data__0__anchor__in,
	input branch_15__phi_n10__valid__0__anchor__in,
	input branch_17__phi_41__ready__0__anchor__in,
	input shl_43__add_44__ready__0__anchor__in,
	input branch_24__Buffer_17__valid__0__anchor__in,
	input cst_18__branch_34__data__0__anchor__in,
	input branchC_55__Buffer_7__data__0__anchor__in,
	input load_80__branch_36__valid__0__anchor__in,
	input fork_0__add_5__valid__0__anchor__in,
	input fork_34__branch_19__ready__0__anchor__in,
	input mul_52__add_53__valid__0__anchor__in,
	input fork_62__phi_42__valid__0__anchor__in,
	input cst_25__MC_A__valid__0__anchor__in,
	input forkC_55__cst_19__valid__0__anchor__in,
	input branch_0__phi_1__ready__0__anchor__in,
	input [31 : 0] z_din0,
	input Buffer_16__phiC_28__ready__0__anchor__in,
	input fork_33__branch_15__valid__0__anchor__in,
	input Buffer_9__phi_36__ready__0__anchor__in,
	input fork_36__branch_29__data__0__anchor__in,
	input brCst_block2__fork_30__ready__0__anchor__in,
	input branch_1__sink_1__valid__0__anchor__in,
	input branch_7__sink_7__ready__0__anchor__in,
	input branch_3__sink_3__data__0__anchor__in,
	input [5 : 0] phi_n13__fork_20__data__0__anchor__in,
	input load_88__mul_89__valid__0__anchor__in,
	input [10 : 0] cst_10__shl_43__data__0__anchor__in,
	input [5 : 0] fork_1__branch_7__data__0__anchor__in,
	input [5 : 0] load_11__MC_u1__data__0__anchor__in,
	input load_22__mul_23__ready__0__anchor__in,
	input branchC_58__phiC_40__ready__0__anchor__in,
	input [31 : 0] branch_12__Buffer_1__data__0__anchor__in,
	input [5 : 0] branch_28__Buffer_9__data__0__anchor__in,
	input fork_37__branch_30__ready__0__anchor__in,
	input fork_36__branch_28__data__0__anchor__in,
	input branch_30__phi_63__valid__0__anchor__in,
	input [31 : 0] phi_n7__branch_10__data__0__anchor__in,
	input fork_62__phi_41__data__0__anchor__in,
	input [5 : 0] fork_9__branch_32__data__0__anchor__in,
	input Buffer_15__phi_n26__ready__0__anchor__in,
	input [31 : 0] branch_1__phi_n0__data__0__anchor__in,
	input fork_31__branch_9__valid__0__anchor__in,
	input fork_35__branch_22__ready__0__anchor__in,
	input branch_3__phi_3__valid__0__anchor__in,
	input [5 : 0] cst_22__icmp_96__data__0__anchor__in,
	input branch_10__Buffer_5__ready__0__anchor__in,
	input load_92__mul_93__valid__0__anchor__in,
	input phiC_40__forkC_57__data__0__anchor__in,
	input phiC_40__forkC_57__valid__0__anchor__in,
	input fork_35__branch_25__ready__0__anchor__in,
	input load_22__mul_23__valid__0__anchor__in,
	input [5 : 0] branch_32__sink_22__data__0__anchor__in,
	input MC_A__load_8__valid__0__anchor__in,
	input branch_31__phi_n20__valid__0__anchor__in,
	input fork_29__branch_0__valid__0__anchor__in,
	input phi_n4__branch_13__ready__0__anchor__in,
	input branch_12__Buffer_1__ready__0__anchor__in,
	input phi_n0__branch_5__ready__0__anchor__in,
	input MC_A__load_8__ready__0__anchor__in,
	input branch_38__sink_27__valid__0__anchor__in,
	input [31 : 0] Buffer_18__phi_n18__data__0__anchor__in,
	input forkC_44__brCst_block1__ready__0__anchor__in,
	input cst_4__add_29__ready__0__anchor__in,
	input phi_n19__branch_31__valid__0__anchor__in,
	input fork_32__branch_11__data__0__anchor__in,
	input MC_x__load_66__valid__0__anchor__in,
	input fork_32__branch_13__valid__0__anchor__in,
	input fork_41__branch_40__data__0__anchor__in,
	input phi_n0__branch_5__valid__0__anchor__in,
	input [31 : 0] load_69__add_70__data__0__anchor__in,
	input fork_62__phi_41__ready__0__anchor__in,
	input branchC_50__phiC_32__ready__0__anchor__in,
	input branchC_59__phiC_41__data__0__anchor__in,
	input branch_12__phi_n8__ready__0__anchor__in,
	input icmp_60__fork_36__data__0__anchor__in,
	input phi_n8__branch_15__valid__0__anchor__in,
	input Buffer_8__phi_82__valid__0__anchor__in,
	input fork_36__branch_27__valid__0__anchor__in,
	input forkC_45__branchC_47__ready__0__anchor__in,
	input [31 : 0] branch_10__phi_n4__data__0__anchor__in,
	input [5 : 0] branch_41__Buffer_29__data__0__anchor__in,
	input branch_16__phi_n11__ready__0__anchor__in,
	input branch_13__phi_n9__ready__0__anchor__in,
	input forkC_55__cst_19__ready__0__anchor__in,
	input [31 : 0] u1_din0,
	input [31 : 0] branch_27__sink_18__data__0__anchor__in,
	input fork_31__branchC_48__data__0__anchor__in,
	input [31 : 0] branch_35__phi_n22__data__0__anchor__in,
	input fork_33__branch_16__ready__0__anchor__in,
	input fork_34__branch_17__valid__0__anchor__in,
	input phiC_29__forkC_46__data__0__anchor__in,
	input fork_40__branchC_57__data__0__anchor__in,
	input MC_y__end_0__data__0__anchor__in,
	input Buffer_23__phi_n27__ready__0__anchor__in,
	input fork_32__branch_12__data__0__anchor__in,
	input [31 : 0] Buffer_1__phi_n0__data__0__anchor__in,
	input branch_23__Buffer_3__ready__0__anchor__in,
	input fork_11__add_95__ready__0__anchor__in,
	input fork_41__branch_42__ready__0__anchor__in,
	input [5 : 0] fork_13__branch_41__data__0__anchor__in,
	input Buffer_6__phiC_38__valid__0__anchor__in,
	input [5 : 0] cst_11__add_54__data__0__anchor__in,
	input icmp_60__fork_36__ready__0__anchor__in,
	input [2 : 0] source_6__cst_10__data__0__anchor__in,
	input phiC_36__forkC_53__ready__0__anchor__in,
	input add_73__fork_9__valid__0__anchor__in,
	input cst_12__icmp_55__ready__0__anchor__in,
	input branch_37__sink_26__valid__0__anchor__in,
	input phi_1__branch_4__valid__0__anchor__in,
	input fork_33__branchC_50__ready__0__anchor__in,
	input branch_15__sink_10__valid__0__anchor__in,
	input Buffer_26__phi_1__valid__0__anchor__in,
	input [31 : 0] branch_43__Buffer_23__data__0__anchor__in,
	input source_12__cst_17__valid__0__anchor__in,
	input fork_38__branch_32__data__0__anchor__in,
	input [5 : 0] add_32__fork_2__data__0__anchor__in,
	input MC_A__load_88__ready__0__anchor__in,
	input [31 : 0] branch_17__phi_41__data__0__anchor__in,
	input phi_41__add_53__ready__0__anchor__in,
	input start_valid,
	input fork_42__branchC_59__valid__0__anchor__in,
	input branch_42__Buffer_15__ready__0__anchor__in,
	input [31 : 0] phi_n6__branch_9__data__0__anchor__in,
	input [5 : 0] load_22__MC_v2__data__0__anchor__in,
	input branch_17__sink_12__ready__0__anchor__in,
	input cst_20__shl_84__valid__0__anchor__in,
	input [5 : 0] fork_0__load_22__data__0__anchor__in,
	input phi_n25__branch_44__ready__0__anchor__in,
	input branchC_56__sink_37__data__0__anchor__in,
	input branchC_53__phiC_35__data__0__anchor__in,
	input source_16__cst_23__valid__0__anchor__in,
	input forkC_44__branchC_46__ready__0__anchor__in,
	input fork_4__shl_43__valid__0__anchor__in,
	input fork_35__branch_24__data__0__anchor__in,
	input branchC_50__sink_34__ready__0__anchor__in,
	input branch_28__sink_19__ready__0__anchor__in,
	input forkC_52__brCst_block9__valid__0__anchor__in,
	input [31 : 0] branch_9__Buffer_4__data__0__anchor__in,
	input branch_10__Buffer_5__valid__0__anchor__in,
	input source_2__cst_4__valid__0__anchor__in,
	input [31 : 0] Buffer_11__phi_n22__data__0__anchor__in,
	input cst_10__shl_43__valid__0__anchor__in,
	input Buffer_17__phi_n16__valid__0__anchor__in,
	input load_92__MC_x__ready__0__anchor__in,
	input [31 : 0] MC_u2__load_19__data__0__anchor__in,
	input fork_31__branch_9__ready__0__anchor__in,
	input forkC_49__brCst_block6__ready__0__anchor__in,
	input icmp_74__fork_38__data__0__anchor__in,
	input Buffer_9__phi_36__valid__0__anchor__in,
	input [5 : 0] branch_3__phi_3__data__0__anchor__in,
	input branch_18__sink_13__data__0__anchor__in,
	input cst_2__shl_4__valid__0__anchor__in,
	input [31 : 0] store_2__MC_x__data__0__anchor__in,
	input fork_0__add_29__ready__0__anchor__in,
	input cst_19__branch_37__data__0__anchor__in,
	input branch_34__sink_23__data__0__anchor__in,
	input forkC_49__cst_9__ready__0__anchor__in,
	input store_1__MC_x__valid__1__anchor__in,
	input Buffer_4__phi_n6__ready__0__anchor__in,
	input add_16__add_24__ready__0__anchor__in,
	input fork_3__branch_21__ready__0__anchor__in,
	input fork_40__branchC_57__valid__0__anchor__in,
	input branch_35__phi_n22__ready__0__anchor__in,
	input branch_14__sink_9__ready__0__anchor__in,
	input [5 : 0] phi_36__fork_3__data__0__anchor__in,
	input branchC_59__Buffer_6__data__0__anchor__in,
	input Buffer_14__phi_n5__ready__0__anchor__in,
	input phi_n6__branch_9__valid__0__anchor__in,
	input cst_4__add_29__valid__0__anchor__in,
	input load_88__MC_A__valid__0__anchor__in,
	input branch_5__phi_n6__valid__0__anchor__in,
	input branch_10__phi_n4__ready__0__anchor__in,
	input [5 : 0] fork_2__icmp_33__data__0__anchor__in,
	input [5 : 0] cst_14__icmp_60__data__0__anchor__in,
	input branch_37__phi_83__valid__0__anchor__in,
	input [31 : 0] branch_16__sink_11__data__0__anchor__in,
	input cst_3__shl_25__valid__0__anchor__in,
	input MC_z__load_69__valid__0__anchor__in,
	input branchC_49__Buffer_16__ready__0__anchor__in,
	input cst_18__branch_34__ready__0__anchor__in,
	input fork_34__branch_19__valid__0__anchor__in,
	input source_14__cst_21__data__0__anchor__in,
	input [31 : 0] load_22__mul_23__data__0__anchor__in,
	input fork_31__branch_7__ready__0__anchor__in,
	input Buffer_28__phi_n20__ready__0__anchor__in,
	input fork_8__add_73__ready__0__anchor__in,
	input cst_13__add_59__valid__0__anchor__in,
	input shl_84__add_85__ready__0__anchor__in,
	input branchC_57__phiC_39__valid__0__anchor__in,
	input Buffer_25__phi_3__valid__0__anchor__in,
	input fork_38__branchC_55__data__0__anchor__in,
	input forkC_52__branchC_54__ready__0__anchor__in,
	input source_0__cst_2__ready__0__anchor__in,
	input fork_42__branch_44__data__0__anchor__in,
	input source_14__cst_21__ready__0__anchor__in,
	input MC_x__load_92__ready__0__anchor__in,
	input [5 : 0] load_66__MC_x__data__0__anchor__in,
	input fork_10__load_80__valid__0__anchor__in,
	input source_8__cst_12__valid__0__anchor__in,
	input branchC_48__phiC_30__valid__0__anchor__in,
	input branch_23__sink_17__ready__0__anchor__in,
	input [5 : 0] fork_11__add_95__data__0__anchor__in,
	input forkC_52__brCst_block9__ready__0__anchor__in,
	input source_15__cst_22__valid__0__anchor__in,
	input fork_38__branch_32__ready__0__anchor__in,
	input add_29__fork_1__ready__0__anchor__in,
	input add_5__load_8__valid__0__anchor__in,
	input [31 : 0] branch_20__phi_n18__data__0__anchor__in,
	input icmp_33__fork_32__valid__0__anchor__in,
	input fork_32__branch_13__ready__0__anchor__in,
	input shl_25__add_26__valid__0__anchor__in,
	input branchC_47__sink_33__data__0__anchor__in,
	input phi_n2__add_32__ready__0__anchor__in,
	input [5 : 0] fork_17__load_11__data__0__anchor__in,
	input branchC_46__sink_32__data__0__anchor__in,
	input [5 : 0] source_15__cst_22__data__0__anchor__in,
	input branchC_53__Buffer_27__ready__0__anchor__in,
	input MC_u2__load_19__valid__0__anchor__in,
	input brCst_block5__fork_33__data__0__anchor__in,
	input [31 : 0] load_51__mul_52__data__0__anchor__in,
	input load_51__mul_52__ready__0__anchor__in,
	input rst,
	input branchC_56__sink_37__valid__0__anchor__in,
	input load_8__add_16__valid__0__anchor__in,
	input fork_30__branch_3__data__0__anchor__in,
	input branchC_53__Buffer_27__data__0__anchor__in,
	input Buffer_18__phi_n18__ready__0__anchor__in,
	input branch_43__phi_n25__valid__0__anchor__in,
	input phi_82__add_94__ready__0__anchor__in,
	input MC_w__end_0__ready__0__anchor__in,
	input shl_43__add_44__valid__0__anchor__in,
	input branch_44__sink_30__valid__0__anchor__in,
	input cst_0__branch_0__valid__0__anchor__in,
	input [31 : 0] phi_n8__branch_15__data__0__anchor__in,
	input [5 : 0] fork_0__add_29__data__0__anchor__in,
	input [31 : 0] MC_A__load_88__data__0__anchor__in,
	input forkC_57__cst_28__data__0__anchor__in,
	input fork_27__branch_42__ready__0__anchor__in,
	input [5 : 0] Buffer_17__phi_n16__data__0__anchor__in,
	input [5 : 0] load_69__MC_z__data__0__anchor__in,
	input branch_23__sink_17__valid__0__anchor__in,
	input fork_29__branchC_46__valid__0__anchor__in,
	input source_6__cst_10__valid__0__anchor__in,
	input phi_36__fork_3__ready__0__anchor__in,
	input [5 : 0] branch_21__sink_16__data__0__anchor__in,
	input [31 : 0] cst_26__MC_x__data__0__anchor__in,
	input [31 : 0] phi_n15__branch_29__data__0__anchor__in,
	input fork_0__load_22__ready__0__anchor__in,
	input branch_40__phi_n23__ready__0__anchor__in,
	input load_39__branch_17__ready__0__anchor__in,
	input phi_3__fork_0__ready__0__anchor__in,
	input phi_n19__branch_31__ready__0__anchor__in,
	input fork_20__add_59__valid__0__anchor__in,
	input forkC_57__branchC_59__valid__0__anchor__in,
	input fork_10__branch_39__valid__0__anchor__in,
	input branch_37__sink_26__data__0__anchor__in,
	input add_53__branch_22__valid__0__anchor__in,
	input fork_31__branch_7__data__0__anchor__in,
	input branchC_59__phiC_41__ready__0__anchor__in,
	input phiC_28__forkC_45__ready__0__anchor__in,
	input branch_9__phi_n3__valid__0__anchor__in,
	input Buffer_10__phi_63__valid__0__anchor__in,
	input add_94__branch_40__valid__0__anchor__in,
	input fork_39__branchC_56__data__0__anchor__in,
	input phi_n5__fork_17__ready__0__anchor__in,
	input add_85__load_88__valid__0__anchor__in,
	input [11 : 0] add_26__store_0__data__0__anchor__in,
	input fork_29__branch_1__ready__0__anchor__in,
	input [5 : 0] phi_83__fork_11__data__0__anchor__in,
	input [5 : 0] source_10__cst_14__data__0__anchor__in,
	input fork_27__shl_84__ready__0__anchor__in,
	input phiC_34__forkC_51__valid__0__anchor__in,
	input branch_37__sink_26__ready__0__anchor__in,
	input [31 : 0] branch_31__sink_21__data__0__anchor__in,
	input MC_w__load_80__ready__0__anchor__in,
	input load_51__MC_y__valid__0__anchor__in,
	input [31 : 0] branch_1__sink_1__data__0__anchor__in,
	input [5 : 0] source_17__cst_24__data__0__anchor__in,
	input [31 : 0] branch_12__phi_n8__data__0__anchor__in,
	input fork_34__branch_20__valid__0__anchor__in,
	input fork_35__branch_24__ready__0__anchor__in,
	input [5 : 0] fork_10__load_80__data__0__anchor__in,
	input icmp_55__fork_35__valid__0__anchor__in,
	input [5 : 0] branch_45__Buffer_0__data__0__anchor__in,
	input store_0__MC_A__valid__0__anchor__in,
	input [31 : 0] load_39__branch_17__data__0__anchor__in,
	input branchC_59__Buffer_6__valid__0__anchor__in,
	input load_11__MC_u1__valid__0__anchor__in,
	input fork_26__store_3__valid__0__anchor__in,
	input phiC_31__forkC_48__ready__0__anchor__in,
	input [11 : 0] add_5__load_8__data__0__anchor__in,
	input load_47__MC_A__ready__0__anchor__in,
	input [31 : 0] load_88__mul_89__data__0__anchor__in,
	input [10 : 0] fork_17__shl_4__data__0__anchor__in,
	input phiC_36__phi_63__valid__0__anchor__in,
	input add_54__fork_6__ready__0__anchor__in,
	input branchC_58__phiC_40__valid__0__anchor__in,
	input fork_6__icmp_55__valid__0__anchor__in,
	input branch_13__Buffer_19__ready__0__anchor__in,
	input branch_19__sink_14__ready__0__anchor__in,
	input cst_24__icmp_101__ready__0__anchor__in,
	input branch_15__phi_n10__ready__0__anchor__in,
	input shl_84__add_85__valid__0__anchor__in,
	input [31 : 0] branch_15__sink_10__data__0__anchor__in,
	input phi_n3__branch_12__valid__0__anchor__in,
	input forkC_55__brCst_block12__ready__0__anchor__in,
	input fork_32__branchC_49__valid__0__anchor__in,
	input fork_11__add_85__ready__0__anchor__in,
	input [5 : 0] branch_34__phi_77__data__0__anchor__in,
	input forkC_54__branchC_56__valid__0__anchor__in,
	input fork_29__branch_0__ready__0__anchor__in,
	input [31 : 0] v2_din1,
	input branch_25__phi_n14__valid__0__anchor__in,
	input cst_16__add_73__ready__0__anchor__in,
	input phiC_37__forkC_54__valid__0__anchor__in,
	input [11 : 0] fork_0__add_5__data__0__anchor__in,
	input [31 : 0] phi_n14__branch_27__data__0__anchor__in,
	input fork_29__branch_2__ready__0__anchor__in,
	input fork_36__branch_27__ready__0__anchor__in,
	input store_2__MC_x__valid__1__anchor__in,
	input [5 : 0] branch_41__sink_29__data__0__anchor__in,
	input fork_41__branch_41__valid__0__anchor__in,
	input cst_9__branch_18__valid__0__anchor__in,
	input [31 : 0] branch_29__phi_n19__data__0__anchor__in,
	input Buffer_13__phi_n10__ready__0__anchor__in,
	input branch_40__phi_n23__valid__0__anchor__in,
	input phi_n14__branch_27__valid__0__anchor__in,
	input [31 : 0] branch_38__sink_27__data__0__anchor__in,
	input forkC_52__cst_15__ready__0__anchor__in,
	input branch_38__phi_n27__ready__0__anchor__in,
	input phi_n11__branch_20__valid__0__anchor__in,
	input [31 : 0] Buffer_8__phi_82__data__0__anchor__in,
	input fork_36__branchC_53__ready__0__anchor__in,
	input cst_16__add_73__valid__0__anchor__in,
	input [31 : 0] phi_n1__branch_6__data__0__anchor__in,
	input branch_2__phi_n1__ready__0__anchor__in,
	input forkC_54__brCst_block11__valid__0__anchor__in,
	input branch_6__sink_6__valid__0__anchor__in,
	input branch_42__Buffer_15__valid__0__anchor__in,
	input forkC_51__branchC_53__ready__0__anchor__in,
	input fork_22__branch_24__valid__0__anchor__in,
	input branch_3__sink_3__ready__0__anchor__in,
	input fork_35__branch_23__valid__0__anchor__in,
	input cst_15__branch_30__ready__0__anchor__in,
	input [31 : 0] add_24__store_0__data__0__anchor__in,
	input [31 : 0] w_din0,
	input branchC_54__sink_36__data__0__anchor__in,
	input Buffer_1__phi_n0__ready__0__anchor__in,
	input fork_30__branchC_47__data__0__anchor__in,
	input fork_1__branch_7__valid__0__anchor__in,
	input [31 : 0] branch_19__sink_14__data__0__anchor__in,
	input fork_28__branch_43__valid__0__anchor__in,
	input cst_0__branch_0__data__0__anchor__in,
	input phi_n27__fork_28__valid__0__anchor__in,
	input branch_30__phi_63__ready__0__anchor__in,
	input forkC_45__cst_1__data__0__anchor__in,
	input forkC_48__branchC_50__data__0__anchor__in,
	input source_8__cst_12__ready__0__anchor__in,
	input branchC_55__Buffer_7__ready__0__anchor__in,
	input branch_28__Buffer_9__valid__0__anchor__in,
	input [31 : 0] MC_x__load_92__data__0__anchor__in,
	input phiC_39__fork_65__valid__0__anchor__in,
	input [31 : 0] MC_x__load_39__data__0__anchor__in,
	input [5 : 0] load_39__MC_x__data__0__anchor__in,
	input branch_29__phi_n19__ready__0__anchor__in,
	input brCst_block6__fork_34__ready__0__anchor__in,
	input forkC_55__branchC_57__data__0__anchor__in,
	input load_80__MC_w__ready__0__anchor__in,
	input branchC_52__phiC_34__valid__0__anchor__in,
	input Buffer_7__phiC_36__ready__0__anchor__in,
	input fork_31__branch_8__data__0__anchor__in,
	input phi_n17__fork_23__valid__0__anchor__in,
	input forkC_49__brCst_block6__valid__0__anchor__in,
	input brCst_block6__fork_34__valid__0__anchor__in,
	input branch_21__phi_n16__valid__0__anchor__in,
	input fork_30__branch_6__valid__0__anchor__in,
	input branch_39__sink_28__valid__0__anchor__in,
	input [5 : 0] fork_20__store_1__data__0__anchor__in,
	input MC_v1__end_0__ready__0__anchor__in,
	input phi_n22__branch_38__valid__0__anchor__in,
	input fork_30__branchC_47__valid__0__anchor__in,
	input [5 : 0] branch_45__sink_31__data__0__anchor__in,
	input [5 : 0] cst_23__add_100__data__0__anchor__in,
	input branch_25__Buffer_22__ready__0__anchor__in,
	input MC_y__end_0__valid__0__anchor__in,
	input [31 : 0] Buffer_5__phi_n7__data__0__anchor__in,
	input add_44__load_47__valid__0__anchor__in,
	input add_59__fork_7__ready__0__anchor__in,
	input cst_17__icmp_74__ready__0__anchor__in,
	input fork_41__branch_43__data__0__anchor__in,
	input alpha_valid_in,
	input [5 : 0] cst_16__add_73__data__0__anchor__in,
	input MC_u1__end_0__valid__0__anchor__in,
	input source_11__cst_16__data__0__anchor__in,
	input [31 : 0] MC_z__load_69__data__0__anchor__in,
	input [5 : 0] phi_n24__fork_26__data__0__anchor__in,
	input add_54__fork_6__valid__0__anchor__in,
	input [5 : 0] branch_0__phi_1__data__0__anchor__in,
	output branchC_46__phiC_28__valid__0__anchor__out,
	output branch_37__sink_26__ready__0__anchor__out,
	output phiC_37__forkC_54__valid__0__anchor__out,
	output [31 : 0] phi_n22__branch_38__data__0__anchor__out,
	output Buffer_11__phi_n22__valid__0__anchor__out,
	output branchC_51__phiC_33__data__0__anchor__out,
	output [31 : 0] branch_2__phi_n1__data__0__anchor__out,
	output phi_n17__fork_23__valid__0__anchor__out,
	output fork_35__branch_24__ready__0__anchor__out,
	output branch_20__sink_15__valid__0__anchor__out,
	output [5 : 0] branch_0__phi_1__data__0__anchor__out,
	output phi_n1__branch_6__ready__0__anchor__out,
	output branchC_50__phiC_32__ready__0__anchor__out,
	output branch_27__Buffer_13__ready__0__anchor__out,
	output [5 : 0] cst_17__icmp_74__data__0__anchor__out,
	output [31 : 0] phi_n1__branch_6__data__0__anchor__out,
	output [5 : 0] fork_7__icmp_60__data__0__anchor__out,
	output branch_12__phi_n8__ready__0__anchor__out,
	output load_80__branch_36__ready__0__anchor__out,
	output phi_n6__branch_9__valid__0__anchor__out,
	output phi_n5__fork_17__valid__0__anchor__out,
	output MC_y__end_0__valid__0__anchor__out,
	output branch_12__phi_n8__valid__0__anchor__out,
	output fork_34__branch_19__ready__0__anchor__out,
	output branch_13__Buffer_19__valid__0__anchor__out,
	output load_66__add_70__valid__0__anchor__out,
	output fork_3__load_39__valid__0__anchor__out,
	output branch_42__phi_n24__valid__0__anchor__out,
	output forkC_48__branchC_50__ready__0__anchor__out,
	output add_24__store_0__ready__0__anchor__out,
	output forkC_57__branchC_59__valid__0__anchor__out,
	output w_ce0,
	output load_22__mul_23__valid__0__anchor__out,
	output phiC_32__forkC_49__ready__0__anchor__out,
	output [31 : 0] phi_n27__fork_28__data__0__anchor__out,
	output icmp_96__fork_41__ready__0__anchor__out,
	output MC_z__load_69__ready__0__anchor__out,
	output [10 : 0] fork_27__shl_84__data__0__anchor__out,
	output fork_17__shl_25__ready__0__anchor__out,
	output cst_9__branch_18__ready__0__anchor__out,
	output forkC_44__branchC_46__data__0__anchor__out,
	output [10 : 0] cst_20__shl_84__data__0__anchor__out,
	output fork_62__phi_41__ready__0__anchor__out,
	output branchC_59__Buffer_6__ready__0__anchor__out,
	output branchC_47__sink_33__valid__0__anchor__out,
	output [31 : 0] phi_n10__branch_19__data__0__anchor__out,
	output [31 : 0] branch_25__phi_n14__data__0__anchor__out,
	output cst_16__add_73__valid__0__anchor__out,
	output phi_n6__branch_9__ready__0__anchor__out,
	output [31 : 0] phi_41__add_53__data__0__anchor__out,
	output forkC_52__cst_15__valid__0__anchor__out,
	output phi_42__fork_4__valid__0__anchor__out,
	output load_11__MC_u1__ready__0__anchor__out,
	output [31 : 0] branch_12__phi_n8__data__0__anchor__out,
	output branch_43__Buffer_23__ready__0__anchor__out,
	output add_53__branch_22__valid__0__anchor__out,
	output phi_n16__fork_22__ready__0__anchor__out,
	output branch_31__phi_n20__ready__0__anchor__out,
	output [5 : 0] phi_36__fork_3__data__0__anchor__out,
	output fork_34__branch_20__ready__0__anchor__out,
	output [5 : 0] store_3__MC_w__data__1__anchor__out,
	output Buffer_7__phiC_36__data__0__anchor__out,
	output load_47__MC_A__valid__0__anchor__out,
	output fork_37__branch_30__data__0__anchor__out,
	output fork_17__load_19__valid__0__anchor__out,
	output load_14__mul_15__valid__0__anchor__out,
	output branchC_49__Buffer_16__data__0__anchor__out,
	output fork_0__add_5__ready__0__anchor__out,
	output [11 : 0] fork_11__add_85__data__0__anchor__out,
	output phi_n7__branch_10__valid__0__anchor__out,
	output MC_A__load_88__ready__0__anchor__out,
	output phiC_30__branchC_49__valid__0__anchor__out,
	output fork_31__branch_7__data__0__anchor__out,
	output MC_x__load_66__ready__0__anchor__out,
	output [31 : 0] x_dout1,
	output [31 : 0] phi_82__add_94__data__0__anchor__out,
	output source_9__cst_13__ready__0__anchor__out,
	output branch_4__phi_n5__valid__0__anchor__out,
	output [5 : 0] fork_27__branch_42__data__0__anchor__out,
	output forkC_49__brCst_block6__data__0__anchor__out,
	output branchC_55__Buffer_7__ready__0__anchor__out,
	output forkC_49__branchC_51__valid__0__anchor__out,
	output fork_29__branch_0__data__0__anchor__out,
	output Buffer_28__phi_n20__valid__0__anchor__out,
	output fork_34__branchC_51__valid__0__anchor__out,
	output Buffer_16__phiC_28__valid__0__anchor__out,
	output start_0__forkC_44__data__0__anchor__out,
	output [11 : 0] store_0__MC_A__data__1__anchor__out,
	output store_2__MC_x__valid__1__anchor__out,
	output mul_93__add_94__valid__0__anchor__out,
	output add_16__add_24__valid__0__anchor__out,
	output branch_35__phi_n22__valid__0__anchor__out,
	output phi_n15__branch_29__ready__0__anchor__out,
	output icmp_74__fork_38__valid__0__anchor__out,
	output [5 : 0] phi_n16__fork_22__data__0__anchor__out,
	output branch_30__sink_20__data__0__anchor__out,
	output cst_2__shl_4__ready__0__anchor__out,
	output [5 : 0] u2_address1,
	output fork_37__branch_31__data__0__anchor__out,
	output branch_32__sink_22__ready__0__anchor__out,
	output Buffer_8__phi_82__valid__0__anchor__out,
	output load_39__branch_17__valid__0__anchor__out,
	output phi_n25__branch_44__ready__0__anchor__out,
	output [11 : 0] A_address1,
	output source_7__cst_11__valid__0__anchor__out,
	output fork_0__load_22__valid__0__anchor__out,
	output cst_25__MC_A__ready__0__anchor__out,
	output x_ce0,
	output branch_43__phi_n25__valid__0__anchor__out,
	output [5 : 0] phi_83__fork_11__data__0__anchor__out,
	output forkC_57__cst_28__valid__0__anchor__out,
	output branchC_48__phiC_30__valid__0__anchor__out,
	output icmp_33__fork_32__valid__0__anchor__out,
	output fork_4__shl_43__ready__0__anchor__out,
	output branch_39__sink_28__valid__0__anchor__out,
	output branch_38__phi_n27__valid__0__anchor__out,
	output branch_8__Buffer_14__valid__0__anchor__out,
	output cst_23__add_100__valid__0__anchor__out,
	output phi_36__fork_3__valid__0__anchor__out,
	output fork_31__branch_10__data__0__anchor__out,
	output fork_1__icmp_30__valid__0__anchor__out,
	output fork_36__branchC_53__valid__0__anchor__out,
	output x_we0,
	output u2_ce0,
	output branch_35__sink_24__valid__0__anchor__out,
	output phi_n2__add_32__ready__0__anchor__out,
	output branch_7__Buffer_25__ready__0__anchor__out,
	output MC_z__end_0__valid__0__anchor__out,
	output fork_17__shl_4__valid__0__anchor__out,
	output phi_n21__branch_35__valid__0__anchor__out,
	output branch_7__Buffer_25__valid__0__anchor__out,
	output [5 : 0] cst_16__add_73__data__0__anchor__out,
	output phi_41__add_53__ready__0__anchor__out,
	output branchC_54__sink_36__data__0__anchor__out,
	output [31 : 0] branch_36__phi_82__data__0__anchor__out,
	output icmp_101__fork_42__data__0__anchor__out,
	output [5 : 0] branch_28__Buffer_9__data__0__anchor__out,
	output [31 : 0] Buffer_22__phi_n17__data__0__anchor__out,
	output fork_23__mul_48__valid__0__anchor__out,
	output branch_18__phi_42__ready__0__anchor__out,
	output [5 : 0] branch_4__phi_n5__data__0__anchor__out,
	output load_8__add_16__valid__0__anchor__out,
	output fork_17__load_11__ready__0__anchor__out,
	output load_92__mul_93__valid__0__anchor__out,
	output load_39__MC_x__valid__0__anchor__out,
	output branchC_54__sink_36__valid__0__anchor__out,
	output branch_15__phi_n10__ready__0__anchor__out,
	output [5 : 0] branch_37__phi_83__data__0__anchor__out,
	output [31 : 0] x_dout0,
	output [31 : 0] branch_43__Buffer_23__data__0__anchor__out,
	output fork_41__branch_41__data__0__anchor__out,
	output fork_29__branchC_46__ready__0__anchor__out,
	output forkC_55__branchC_57__data__0__anchor__out,
	output [31 : 0] branch_10__phi_n4__data__0__anchor__out,
	output phi_82__add_94__valid__0__anchor__out,
	output phiC_30__branchC_49__ready__0__anchor__out,
	output [5 : 0] cst_21__add_95__data__0__anchor__out,
	output [5 : 0] branch_21__phi_n16__data__0__anchor__out,
	output [11 : 0] shl_43__add_44__data__0__anchor__out,
	output fork_33__branch_16__data__0__anchor__out,
	output [11 : 0] add_44__load_47__data__0__anchor__out,
	output fork_29__branch_1__valid__0__anchor__out,
	output fork_42__branchC_59__data__0__anchor__out,
	output branchC_58__phiC_40__valid__0__anchor__out,
	output fork_2__icmp_33__valid__0__anchor__out,
	output branch_4__sink_4__ready__0__anchor__out,
	output fork_35__branch_22__ready__0__anchor__out,
	output branchC_54__sink_36__ready__0__anchor__out,
	output MC_v1__end_0__ready__0__anchor__out,
	output [5 : 0] source_17__cst_24__data__0__anchor__out,
	output y_we1,
	output [5 : 0] store_2__MC_x__data__1__anchor__out,
	output cst_1__branch_3__data__0__anchor__out,
	output branch_34__phi_77__valid__0__anchor__out,
	output MC_v1__load_14__valid__0__anchor__out,
	output [5 : 0] branch_11__Buffer_26__data__0__anchor__out,
	output [31 : 0] branch_27__Buffer_13__data__0__anchor__out,
	output branch_36__sink_25__ready__0__anchor__out,
	output branch_31__sink_21__ready__0__anchor__out,
	output phiC_33__fork_62__ready__0__anchor__out,
	output fork_65__phi_82__data__0__anchor__out,
	output phi_n11__branch_20__valid__0__anchor__out,
	output fork_28__mul_89__valid__0__anchor__out,
	output [31 : 0] branch_2__sink_2__data__0__anchor__out,
	output branch_16__sink_11__ready__0__anchor__out,
	output source_6__cst_10__valid__0__anchor__out,
	output [5 : 0] cst_13__add_59__data__0__anchor__out,
	output source_4__cst_6__ready__0__anchor__out,
	output fork_7__branch_28__ready__0__anchor__out,
	output forkC_54__branchC_56__valid__0__anchor__out,
	output [31 : 0] Buffer_19__phi_n1__data__0__anchor__out,
	output ret_0__end_0__ready__0__anchor__out,
	output [5 : 0] u1_address1,
	output [31 : 0] phi_n8__branch_15__data__0__anchor__out,
	output fork_32__branchC_49__valid__0__anchor__out,
	output [5 : 0] fork_26__add_100__data__0__anchor__out,
	output [31 : 0] branch_9__phi_n3__data__0__anchor__out,
	output cst_7__icmp_33__valid__0__anchor__out,
	output load_80__MC_w__ready__0__anchor__out,
	output phi_n11__branch_20__ready__0__anchor__out,
	output [5 : 0] fork_8__add_73__data__0__anchor__out,
	output fork_34__branch_21__data__0__anchor__out,
	output phi_n1__branch_6__valid__0__anchor__out,
	output fork_31__branch_8__data__0__anchor__out,
	output fork_2__branch_11__ready__0__anchor__out,
	output [31 : 0] MC_y__load_51__data__0__anchor__out,
	output brCst_block9__fork_37__valid__0__anchor__out,
	output [31 : 0] branch_1__phi_n0__data__0__anchor__out,
	output load_66__MC_x__valid__0__anchor__out,
	output [31 : 0] branch_44__Buffer_11__data__0__anchor__out,
	output phiC_36__phi_63__data__0__anchor__out,
	output MC_x__load_92__valid__0__anchor__out,
	output forkC_49__cst_9__valid__0__anchor__out,
	output store_0__MC_A__ready__1__anchor__out,
	output branchC_49__phiC_31__valid__0__anchor__out,
	output Buffer_29__phi_83__valid__0__anchor__out,
	output phiC_39__fork_65__ready__0__anchor__out,
	output branch_0__phi_1__ready__0__anchor__out,
	output MC_y__load_51__valid__0__anchor__out,
	output fork_34__branch_17__valid__0__anchor__out,
	output store_2__MC_x__ready__1__anchor__out,
	output fork_13__icmp_96__ready__0__anchor__out,
	output [31 : 0] MC_z__load_69__data__0__anchor__out,
	output forkC_54__brCst_block11__ready__0__anchor__out,
	output phiC_38__phi_77__valid__0__anchor__out,
	output [31 : 0] Buffer_24__phi_n11__data__0__anchor__out,
	output [5 : 0] v2_address0,
	output brCst_block6__fork_34__ready__0__anchor__out,
	output fork_6__branch_23__ready__0__anchor__out,
	output forkC_53__branchC_55__ready__0__anchor__out,
	output [31 : 0] u1_dout0,
	output [31 : 0] alpha__branch_2__data__0__anchor__out,
	output branch_2__phi_n1__ready__0__anchor__out,
	output branchC_54__phiC_36__ready__0__anchor__out,
	output load_47__mul_48__ready__0__anchor__out,
	output branch_25__phi_n14__valid__0__anchor__out,
	output Buffer_27__phiC_32__valid__0__anchor__out,
	output Buffer_8__phi_82__ready__0__anchor__out,
	output phiC_28__phi_1__ready__0__anchor__out,
	output branch_19__sink_14__ready__0__anchor__out,
	output cst_0__branch_0__valid__0__anchor__out,
	output phi_n14__branch_27__ready__0__anchor__out,
	output fork_8__add_73__valid__0__anchor__out,
	output fork_38__branchC_55__data__0__anchor__out,
	output [31 : 0] branch_16__sink_11__data__0__anchor__out,
	output forkC_44__brCst_block1__valid__0__anchor__out,
	output fork_6__icmp_55__valid__0__anchor__out,
	output Buffer_1__phi_n0__valid__0__anchor__out,
	output source_11__cst_16__data__0__anchor__out,
	output A_we0,
	output [5 : 0] branch_4__sink_4__data__0__anchor__out,
	output fork_40__branch_37__ready__0__anchor__out,
	output cst_17__icmp_74__valid__0__anchor__out,
	output add_94__branch_40__valid__0__anchor__out,
	output fork_30__branch_5__data__0__anchor__out,
	output [5 : 0] fork_1__icmp_30__data__0__anchor__out,
	output [2 : 0] source_6__cst_10__data__0__anchor__out,
	output [5 : 0] z_address0,
	output brCst_block9__fork_37__ready__0__anchor__out,
	output store_3__MC_w__ready__1__anchor__out,
	output branch_25__Buffer_22__valid__0__anchor__out,
	output Buffer_13__phi_n10__ready__0__anchor__out,
	output Buffer_20__phiC_29__valid__0__anchor__out,
	output phi_36__fork_3__ready__0__anchor__out,
	output fork_27__branch_42__ready__0__anchor__out,
	output cst_8__branch_14__ready__0__anchor__out,
	output [5 : 0] Buffer_15__phi_n26__data__0__anchor__out,
	output branch_13__Buffer_19__ready__0__anchor__out,
	output fork_62__phi_41__data__0__anchor__out,
	output fork_8__store_2__ready__0__anchor__out,
	output forkC_49__brCst_block6__valid__0__anchor__out,
	output branchC_52__Buffer_21__ready__0__anchor__out,
	output [5 : 0] Buffer_14__phi_n5__data__0__anchor__out,
	output forkC_54__brCst_block11__data__0__anchor__out,
	output branch_11__Buffer_26__valid__0__anchor__out,
	output [5 : 0] branch_14__phi_36__data__0__anchor__out,
	output fork_39__branch_34__data__0__anchor__out,
	output [31 : 0] fork_23__branch_25__data__0__anchor__out,
	output branch_15__sink_10__ready__0__anchor__out,
	output fork_33__branch_14__ready__0__anchor__out,
	output phiC_33__fork_62__valid__0__anchor__out,
	output source_17__cst_24__ready__0__anchor__out,
	output branch_29__Buffer_24__ready__0__anchor__out,
	output Buffer_7__phiC_36__valid__0__anchor__out,
	output shl_25__add_26__ready__0__anchor__out,
	output [31 : 0] phi_n20__branch_33__data__0__anchor__out,
	output add_24__store_0__valid__0__anchor__out,
	output fork_62__phi_42__ready__0__anchor__out,
	output branch_37__sink_26__data__0__anchor__out,
	output fork_29__branch_1__ready__0__anchor__out,
	output forkC_46__cst_25__data__0__anchor__out,
	output add_5__load_8__valid__0__anchor__out,
	output phi_n7__branch_10__ready__0__anchor__out,
	output [31 : 0] y_dout1,
	output branch_3__sink_3__valid__0__anchor__out,
	output fork_26__store_3__ready__0__anchor__out,
	output phi_n10__branch_19__ready__0__anchor__out,
	output phi_83__fork_11__ready__0__anchor__out,
	output [5 : 0] branch_21__sink_16__data__0__anchor__out,
	output load_39__branch_17__ready__0__anchor__out,
	output [5 : 0] phi_n13__fork_20__data__0__anchor__out,
	output shl_43__add_44__valid__0__anchor__out,
	output branch_33__phi_n21__valid__0__anchor__out,
	output [5 : 0] fork_3__branch_21__data__0__anchor__out,
	output Buffer_13__phi_n10__valid__0__anchor__out,
	output fork_34__branch_19__data__0__anchor__out,
	output phiC_39__fork_65__valid__0__anchor__out,
	output forkC_44__cst_0__valid__0__anchor__out,
	output fork_8__load_69__valid__0__anchor__out,
	output [5 : 0] fork_10__branch_39__data__0__anchor__out,
	output branchC_46__sink_32__ready__0__anchor__out,
	output cst_24__icmp_101__ready__0__anchor__out,
	output mul_15__add_16__valid__0__anchor__out,
	output MC_u1__end_0__valid__0__anchor__out,
	output phiC_29__forkC_46__valid__0__anchor__out,
	output MC_w__end_0__ready__0__anchor__out,
	output [31 : 0] branch_17__phi_41__data__0__anchor__out,
	output source_16__cst_23__ready__0__anchor__out,
	output add_85__load_88__valid__0__anchor__out,
	output phiC_28__forkC_45__data__0__anchor__out,
	output fork_41__branch_42__valid__0__anchor__out,
	output forkC_51__branchC_53__data__0__anchor__out,
	output phiC_38__Buffer_30__valid__0__anchor__out,
	output fork_27__shl_84__ready__0__anchor__out,
	output start_0__forkC_44__valid__0__anchor__out,
	output branchC_47__phiC_29__valid__0__anchor__out,
	output [31 : 0] branch_31__sink_21__data__0__anchor__out,
	output cst_3__shl_25__ready__0__anchor__out,
	output store_1__MC_x__valid__1__anchor__out,
	output fork_33__branch_14__data__0__anchor__out,
	output u2_we0,
	output branch_4__sink_4__valid__0__anchor__out,
	output forkC_53__cst_27__valid__0__anchor__out,
	output forkC_55__brCst_block12__data__0__anchor__out,
	output [5 : 0] cst_12__icmp_55__data__0__anchor__out,
	output [31 : 0] store_2__MC_x__data__0__anchor__out,
	output [5 : 0] source_15__cst_22__data__0__anchor__out,
	output branch_28__Buffer_9__valid__0__anchor__out,
	output branchC_59__phiC_41__data__0__anchor__out,
	output MC_A__end_0__data__0__anchor__out,
	output add_5__load_8__ready__0__anchor__out,
	output fork_40__branch_37__data__0__anchor__out,
	output source_14__cst_21__ready__0__anchor__out,
	output load_19__mul_23__ready__0__anchor__out,
	output [31 : 0] mul_93__add_94__data__0__anchor__out,
	output phiC_38__Buffer_30__ready__0__anchor__out,
	output branch_9__Buffer_4__valid__0__anchor__out,
	output fork_33__branch_15__data__0__anchor__out,
	output forkC_53__cst_27__ready__0__anchor__out,
	output fork_22__branch_24__ready__0__anchor__out,
	output phiC_41__ret_0__valid__0__anchor__out,
	output fork_30__branch_6__ready__0__anchor__out,
	output [31 : 0] branch_43__phi_n25__data__0__anchor__out,
	output fork_34__branch_17__ready__0__anchor__out,
	output Buffer_14__phi_n5__ready__0__anchor__out,
	output cst_0__branch_0__data__0__anchor__out,
	output fork_32__branch_11__ready__0__anchor__out,
	output [31 : 0] v2_dout0,
	output branch_6__sink_6__valid__0__anchor__out,
	output branch_27__sink_18__ready__0__anchor__out,
	output x_ce1,
	output branch_43__Buffer_23__valid__0__anchor__out,
	output [31 : 0] branch_9__Buffer_4__data__0__anchor__out,
	output branchC_47__phiC_29__ready__0__anchor__out,
	output fork_26__add_100__ready__0__anchor__out,
	output phiC_31__forkC_48__valid__0__anchor__out,
	output phi_n0__branch_5__valid__0__anchor__out,
	output phi_n9__branch_16__ready__0__anchor__out,
	output A_we1,
	output fork_35__branch_25__valid__0__anchor__out,
	output cst_6__add_32__valid__0__anchor__out,
	output branch_17__sink_12__ready__0__anchor__out,
	output [31 : 0] load_80__branch_36__data__0__anchor__out,
	output Buffer_19__phi_n1__valid__0__anchor__out,
	output branchC_53__Buffer_27__ready__0__anchor__out,
	output source_10__cst_14__ready__0__anchor__out,
	output fork_34__branch_20__valid__0__anchor__out,
	output cst_17__icmp_74__ready__0__anchor__out,
	output branch_24__Buffer_17__valid__0__anchor__out,
	output v1_we1,
	output fork_14__branch_45__ready__0__anchor__out,
	output source_12__cst_17__ready__0__anchor__out,
	output cst_19__branch_37__ready__0__anchor__out,
	output branchC_48__Buffer_20__ready__0__anchor__out,
	output source_13__cst_20__valid__0__anchor__out,
	output [31 : 0] branch_15__phi_n10__data__0__anchor__out,
	output branch_15__phi_n10__valid__0__anchor__out,
	output [31 : 0] load_14__mul_15__data__0__anchor__out,
	output branchC_53__phiC_35__valid__0__anchor__out,
	output branch_37__sink_26__valid__0__anchor__out,
	output fork_62__phi_42__valid__0__anchor__out,
	output Buffer_9__phi_36__valid__0__anchor__out,
	output phiC_40__forkC_57__data__0__anchor__out,
	output branchC_57__sink_38__data__0__anchor__out,
	output brCst_block11__fork_39__valid__0__anchor__out,
	output icmp_30__fork_31__valid__0__anchor__out,
	output fork_42__branch_45__ready__0__anchor__out,
	output forkC_45__branchC_47__data__0__anchor__out,
	output forkC_51__branchC_53__valid__0__anchor__out,
	output Buffer_27__phiC_32__data__0__anchor__out,
	output A_ce1,
	output branch_12__Buffer_1__valid__0__anchor__out,
	output phi_n27__fork_28__ready__0__anchor__out,
	output [5 : 0] fork_10__load_80__data__0__anchor__out,
	output fork_30__branch_6__valid__0__anchor__out,
	output phi_n8__branch_15__ready__0__anchor__out,
	output fork_40__branchC_57__ready__0__anchor__out,
	output [5 : 0] load_22__MC_v2__data__0__anchor__out,
	output branch_35__sink_24__ready__0__anchor__out,
	output [31 : 0] phi_n12__store_1__data__0__anchor__out,
	output [5 : 0] cst_23__add_100__data__0__anchor__out,
	output branch_21__phi_n16__ready__0__anchor__out,
	output phi_n27__fork_28__valid__0__anchor__out,
	output Buffer_20__phiC_29__ready__0__anchor__out,
	output Buffer_22__phi_n17__ready__0__anchor__out,
	output [5 : 0] branch_39__phi_n26__data__0__anchor__out,
	output [31 : 0] branch_27__sink_18__data__0__anchor__out,
	output phiC_40__forkC_57__ready__0__anchor__out,
	output load_51__mul_52__ready__0__anchor__out,
	output add_53__branch_22__ready__0__anchor__out,
	output fork_13__icmp_96__valid__0__anchor__out,
	output phi_n22__branch_38__valid__0__anchor__out,
	output Buffer_25__phi_3__ready__0__anchor__out,
	output Buffer_30__forkC_55__ready__0__anchor__out,
	output fork_11__add_85__ready__0__anchor__out,
	output fork_39__branch_34__valid__0__anchor__out,
	output branch_44__Buffer_11__valid__0__anchor__out,
	output phiC_35__forkC_52__data__0__anchor__out,
	output [5 : 0] branch_32__Buffer_10__data__0__anchor__out,
	output cst_27__MC_x__ready__0__anchor__out,
	output load_69__MC_z__ready__0__anchor__out,
	output forkC_54__branchC_56__data__0__anchor__out,
	output fork_35__branch_23__data__0__anchor__out,
	output fork_37__branchC_54__data__0__anchor__out,
	output [31 : 0] Buffer_4__phi_n6__data__0__anchor__out,
	output cst_15__branch_30__valid__0__anchor__out,
	output branch_41__Buffer_29__ready__0__anchor__out,
	output branch_14__sink_9__ready__0__anchor__out,
	output store_2__MC_x__valid__0__anchor__out,
	output forkC_49__cst_9__data__0__anchor__out,
	output [5 : 0] branch_42__Buffer_15__data__0__anchor__out,
	output branch_16__phi_n11__ready__0__anchor__out,
	output [5 : 0] branch_28__sink_19__data__0__anchor__out,
	output fork_31__branchC_48__valid__0__anchor__out,
	output icmp_60__fork_36__data__0__anchor__out,
	output cst_14__icmp_60__valid__0__anchor__out,
	output store_1__MC_x__ready__0__anchor__out,
	output fork_29__branch_2__ready__0__anchor__out,
	output branch_26__Buffer_18__ready__0__anchor__out,
	output [31 : 0] MC_A__load_47__data__0__anchor__out,
	output fork_38__branch_32__ready__0__anchor__out,
	output fork_40__branch_38__valid__0__anchor__out,
	output phi_n0__branch_5__ready__0__anchor__out,
	output forkC_44__brCst_block1__ready__0__anchor__out,
	output [5 : 0] cst_14__icmp_60__data__0__anchor__out,
	output branchC_49__Buffer_16__ready__0__anchor__out,
	output icmp_55__fork_35__ready__0__anchor__out,
	output phi_n18__branch_26__ready__0__anchor__out,
	output fork_33__branchC_50__data__0__anchor__out,
	output brCst_block12__fork_40__ready__0__anchor__out,
	output [10 : 0] cst_10__shl_43__data__0__anchor__out,
	output [5 : 0] store_1__MC_x__data__1__anchor__out,
	output branch_33__Buffer_28__ready__0__anchor__out,
	output branch_26__phi_n15__valid__0__anchor__out,
	output shl_43__add_44__ready__0__anchor__out,
	output fork_10__load_80__ready__0__anchor__out,
	output branch_45__sink_31__valid__0__anchor__out,
	output forkC_45__cst_1__ready__0__anchor__out,
	output fork_34__branch_18__valid__0__anchor__out,
	output phiC_31__forkC_48__ready__0__anchor__out,
	output [5 : 0] fork_2__branch_11__data__0__anchor__out,
	output fork_41__branch_43__ready__0__anchor__out,
	output [5 : 0] v1_address0,
	output z_we1,
	output fork_38__branch_33__data__0__anchor__out,
	output [5 : 0] x_address0,
	output branch_14__sink_9__valid__0__anchor__out,
	output [31 : 0] branch_5__sink_5__data__0__anchor__out,
	output [11 : 0] load_47__MC_A__data__0__anchor__out,
	output [31 : 0] branch_16__phi_n11__data__0__anchor__out,
	output cst_9__branch_18__data__0__anchor__out,
	output forkC_52__branchC_54__ready__0__anchor__out,
	output branch_5__sink_5__ready__0__anchor__out,
	output source_5__cst_7__valid__0__anchor__out,
	output branch_6__phi_n7__ready__0__anchor__out,
	output fork_42__branchC_59__valid__0__anchor__out,
	output branch_39__phi_n26__valid__0__anchor__out,
	output fork_4__add_54__ready__0__anchor__out,
	output Buffer_10__phi_63__valid__0__anchor__out,
	output brCst_block5__fork_33__data__0__anchor__out,
	output fork_17__shl_25__valid__0__anchor__out,
	output fork_10__branch_39__ready__0__anchor__out,
	output fork_40__branch_36__valid__0__anchor__out,
	output forkC_48__brCst_block5__ready__0__anchor__out,
	output [31 : 0] Buffer_30__forkC_55__data__0__anchor__out,
	output MC_v2__end_0__valid__0__anchor__out,
	output forkC_55__cst_19__ready__0__anchor__out,
	output branch_14__sink_9__data__0__anchor__out,
	output forkC_48__brCst_block5__data__0__anchor__out,
	output Buffer_25__phi_3__valid__0__anchor__out,
	output branch_9__phi_n3__ready__0__anchor__out,
	output fork_36__branch_28__data__0__anchor__out,
	output icmp_55__fork_35__valid__0__anchor__out,
	output fork_4__load_51__ready__0__anchor__out,
	output MC_z__end_0__data__0__anchor__out,
	output [5 : 0] fork_17__branch_8__data__0__anchor__out,
	output Buffer_27__phiC_32__ready__0__anchor__out,
	output fork_30__branch_3__valid__0__anchor__out,
	output branchC_48__Buffer_20__valid__0__anchor__out,
	output [31 : 0] branch_35__phi_n22__data__0__anchor__out,
	output branchC_51__sink_35__ready__0__anchor__out,
	output MC_u2__load_19__valid__0__anchor__out,
	output branch_5__phi_n6__valid__0__anchor__out,
	output [11 : 0] shl_4__add_5__data__0__anchor__out,
	output fork_31__branch_10__valid__0__anchor__out,
	output source_4__cst_6__valid__0__anchor__out,
	output fork_28__mul_89__ready__0__anchor__out,
	output fork_30__branchC_47__ready__0__anchor__out,
	output fork_28__branch_43__ready__0__anchor__out,
	output fork_35__branch_22__valid__0__anchor__out,
	output fork_34__branchC_51__ready__0__anchor__out,
	output branch_6__sink_6__ready__0__anchor__out,
	output fork_39__branchC_56__valid__0__anchor__out,
	output MC_w__load_80__valid__0__anchor__out,
	output fork_34__branch_18__data__0__anchor__out,
	output forkC_46__cst_25__valid__0__anchor__out,
	output MC_v1__load_14__ready__0__anchor__out,
	output store_1__MC_x__ready__1__anchor__out,
	output load_51__MC_y__ready__0__anchor__out,
	output MC_x__load_39__valid__0__anchor__out,
	output forkC_48__cst_8__valid__0__anchor__out,
	output MC_v2__load_22__ready__0__anchor__out,
	output forkC_45__brCst_block2__ready__0__anchor__out,
	output [31 : 0] mul_15__add_16__data__0__anchor__out,
	output branchC_57__phiC_39__data__0__anchor__out,
	output source_5__cst_7__ready__0__anchor__out,
	output MC_z__load_69__valid__0__anchor__out,
	output branch_36__sink_25__valid__0__anchor__out,
	output [31 : 0] cst_28__MC_w__data__0__anchor__out,
	output MC_u1__end_0__data__0__anchor__out,
	output Buffer_23__phi_n27__valid__0__anchor__out,
	output phiC_35__forkC_52__valid__0__anchor__out,
	output [31 : 0] phi_n25__branch_44__data__0__anchor__out,
	output [31 : 0] branch_38__sink_27__data__0__anchor__out,
	output add_54__fork_6__valid__0__anchor__out,
	output [31 : 0] load_92__mul_93__data__0__anchor__out,
	output branch_2__phi_n1__valid__0__anchor__out,
	output fork_65__phi_82__valid__0__anchor__out,
	output phi_63__fork_8__valid__0__anchor__out,
	output branch_41__sink_29__valid__0__anchor__out,
	output branch_35__phi_n22__ready__0__anchor__out,
	output phiC_35__forkC_52__ready__0__anchor__out,
	output [5 : 0] fork_9__branch_32__data__0__anchor__out,
	output mul_23__add_24__valid__0__anchor__out,
	output [31 : 0] branch_19__sink_14__data__0__anchor__out,
	output [31 : 0] MC_x__load_92__data__0__anchor__out,
	output fork_37__branch_30__ready__0__anchor__out,
	output fork_39__branchC_56__ready__0__anchor__out,
	output load_69__add_70__ready__0__anchor__out,
	output [5 : 0] source_8__cst_12__data__0__anchor__out,
	output [5 : 0] fork_11__add_95__data__0__anchor__out,
	output branch_22__phi_n12__ready__0__anchor__out,
	output MC_A__load_8__ready__0__anchor__out,
	output fork_31__branch_7__valid__0__anchor__out,
	output fork_35__branch_23__valid__0__anchor__out,
	output [11 : 0] add_85__load_88__data__0__anchor__out,
	output fork_11__add_95__ready__0__anchor__out,
	output add_95__fork_13__valid__0__anchor__out,
	output [5 : 0] cst_22__icmp_96__data__0__anchor__out,
	output [5 : 0] branch_39__sink_28__data__0__anchor__out,
	output forkC_53__branchC_55__valid__0__anchor__out,
	output Buffer_9__phi_36__ready__0__anchor__out,
	output branch_40__Buffer_8__valid__0__anchor__out,
	output [5 : 0] source_10__cst_14__data__0__anchor__out,
	output branchC_52__phiC_34__data__0__anchor__out,
	output fork_42__branch_44__ready__0__anchor__out,
	output [31 : 0] cst_26__MC_x__data__0__anchor__out,
	output branch_9__Buffer_4__ready__0__anchor__out,
	output phiC_29__forkC_46__data__0__anchor__out,
	output branchC_51__phiC_33__ready__0__anchor__out,
	output branch_18__sink_13__valid__0__anchor__out,
	output cst_15__branch_30__data__0__anchor__out,
	output branchC_52__Buffer_21__valid__0__anchor__out,
	output add_94__branch_40__ready__0__anchor__out,
	output source_1__cst_3__ready__0__anchor__out,
	output cst_13__add_59__ready__0__anchor__out,
	output MC_y__end_0__ready__0__anchor__out,
	output cst_3__shl_25__valid__0__anchor__out,
	output MC_A__load_47__valid__0__anchor__out,
	output cst_25__MC_A__valid__0__anchor__out,
	output fork_8__store_2__valid__0__anchor__out,
	output fork_33__branch_15__ready__0__anchor__out,
	output branch_1__phi_n0__ready__0__anchor__out,
	output branch_20__sink_15__ready__0__anchor__out,
	output Buffer_5__phi_n7__ready__0__anchor__out,
	output forkC_54__cst_18__data__0__anchor__out,
	output brCst_block2__fork_30__valid__0__anchor__out,
	output fork_65__phi_83__valid__0__anchor__out,
	output fork_65__phi_83__data__0__anchor__out,
	output branch_5__phi_n6__ready__0__anchor__out,
	output [31 : 0] branch_33__Buffer_28__data__0__anchor__out,
	output source_8__cst_12__ready__0__anchor__out,
	output [31 : 0] Buffer_23__phi_n27__data__0__anchor__out,
	output branch_17__phi_41__valid__0__anchor__out,
	output add_26__store_0__valid__0__anchor__out,
	output branchC_52__Buffer_21__data__0__anchor__out,
	output forkC_57__cst_28__data__0__anchor__out,
	output [5 : 0] phi_3__fork_0__data__0__anchor__out,
	output [31 : 0] cst_27__MC_x__data__0__anchor__out,
	output forkC_54__cst_18__ready__0__anchor__out,
	output source_2__cst_4__valid__0__anchor__out,
	output [31 : 0] branch_33__phi_n21__data__0__anchor__out,
	output branch_34__sink_23__data__0__anchor__out,
	output [11 : 0] load_88__MC_A__data__0__anchor__out,
	output [5 : 0] fork_13__branch_41__data__0__anchor__out,
	output [31 : 0] branch_6__sink_6__data__0__anchor__out,
	output [5 : 0] load_51__MC_y__data__0__anchor__out,
	output phi_77__fork_10__ready__0__anchor__out,
	output fork_29__branch_1__data__0__anchor__out,
	output forkC_48__cst_8__ready__0__anchor__out,
	output forkC_54__brCst_block11__valid__0__anchor__out,
	output [11 : 0] fork_22__add_44__data__0__anchor__out,
	output load_80__MC_w__valid__0__anchor__out,
	output [5 : 0] fork_17__load_19__data__0__anchor__out,
	output store_1__MC_x__valid__0__anchor__out,
	output [31 : 0] v1_dout0,
	output [31 : 0] branch_29__Buffer_24__data__0__anchor__out,
	output fork_20__add_59__ready__0__anchor__out,
	output [31 : 0] branch_26__phi_n15__data__0__anchor__out,
	output fork_10__load_80__valid__0__anchor__out,
	output [31 : 0] branch_35__sink_24__data__0__anchor__out,
	output phi_n23__store_3__valid__0__anchor__out,
	output brCst_block6__fork_34__valid__0__anchor__out,
	output branchC_54__phiC_36__valid__0__anchor__out,
	output x_we1,
	output [31 : 0] branch_6__phi_n7__data__0__anchor__out,
	output MC_w__load_80__ready__0__anchor__out,
	output [31 : 0] branch_44__sink_30__data__0__anchor__out,
	output fork_42__branch_44__valid__0__anchor__out,
	output phiC_36__forkC_53__ready__0__anchor__out,
	output [5 : 0] fork_14__branch_45__data__0__anchor__out,
	output Buffer_30__forkC_55__valid__0__anchor__out,
	output load_92__MC_x__valid__0__anchor__out,
	output branch_38__phi_n27__ready__0__anchor__out,
	output w_we0,
	output [5 : 0] Buffer_29__phi_83__data__0__anchor__out,
	output [5 : 0] fork_20__store_1__data__0__anchor__out,
	output fork_32__branch_12__data__0__anchor__out,
	output fork_29__branchC_46__data__0__anchor__out,
	output phiC_36__forkC_53__valid__0__anchor__out,
	output [31 : 0] branch_17__sink_12__data__0__anchor__out,
	output [31 : 0] load_47__mul_48__data__0__anchor__out,
	output u2_we1,
	output forkC_44__brCst_block1__data__0__anchor__out,
	output fork_41__branch_42__ready__0__anchor__out,
	output branch_3__sink_3__ready__0__anchor__out,
	output forkC_52__brCst_block9__valid__0__anchor__out,
	output forkC_51__branchC_53__ready__0__anchor__out,
	output [31 : 0] Buffer_28__phi_n20__data__0__anchor__out,
	output [5 : 0] cst_11__add_54__data__0__anchor__out,
	output MC_u1__load_11__ready__0__anchor__out,
	output phiC_36__phi_63__valid__0__anchor__out,
	output fork_35__branch_26__valid__0__anchor__out,
	output forkC_48__branchC_50__valid__0__anchor__out,
	output fork_33__branchC_50__ready__0__anchor__out,
	output branch_2__sink_2__valid__0__anchor__out,
	output v2_ce1,
	output [31 : 0] MC_v1__load_14__data__0__anchor__out,
	output phi_3__fork_0__ready__0__anchor__out,
	output branchC_58__phiC_40__data__0__anchor__out,
	output branch_22__Buffer_12__ready__0__anchor__out,
	output [31 : 0] mul_48__mul_52__data__0__anchor__out,
	output forkC_55__brCst_block12__valid__0__anchor__out,
	output fork_42__branch_45__data__0__anchor__out,
	output fork_34__branch_20__data__0__anchor__out,
	output add_70__store_2__ready__0__anchor__out,
	output [31 : 0] load_66__add_70__data__0__anchor__out,
	output fork_7__branch_28__valid__0__anchor__out,
	output branch_40__phi_n23__ready__0__anchor__out,
	output forkC_46__cst_25__ready__0__anchor__out,
	output [5 : 0] load_69__MC_z__data__0__anchor__out,
	output [31 : 0] phi_n14__branch_27__data__0__anchor__out,
	output source_14__cst_21__valid__0__anchor__out,
	output branch_1__sink_1__valid__0__anchor__out,
	output store_3__MC_w__valid__1__anchor__out,
	output phi_n13__fork_20__ready__0__anchor__out,
	output [5 : 0] fork_4__load_51__data__0__anchor__out,
	output phiC_30__branchC_49__data__0__anchor__out,
	output cst_28__MC_w__valid__0__anchor__out,
	output branch_16__phi_n11__valid__0__anchor__out,
	output fork_62__phi_42__data__0__anchor__out,
	output add_54__fork_6__ready__0__anchor__out,
	output add_26__store_0__ready__0__anchor__out,
	output fork_38__branch_32__data__0__anchor__out,
	output fork_17__branch_8__ready__0__anchor__out,
	output cst_20__shl_84__valid__0__anchor__out,
	output fork_11__load_92__ready__0__anchor__out,
	output [5 : 0] add_32__fork_2__data__0__anchor__out,
	output cst_5__icmp_30__valid__0__anchor__out,
	output fork_13__branch_41__ready__0__anchor__out,
	output source_16__cst_23__valid__0__anchor__out,
	output [11 : 0] fork_0__add_5__data__0__anchor__out,
	output phiC_33__fork_62__data__0__anchor__out,
	output MC_w__end_0__valid__0__anchor__out,
	output MC_z__end_0__ready__0__anchor__out,
	output branchC_59__Buffer_6__valid__0__anchor__out,
	output phi_n15__branch_29__valid__0__anchor__out,
	output branch_18__sink_13__data__0__anchor__out,
	output [11 : 0] shl_84__add_85__data__0__anchor__out,
	output branch_23__Buffer_3__ready__0__anchor__out,
	output [5 : 0] branch_41__sink_29__data__0__anchor__out,
	output Buffer_18__phi_n18__ready__0__anchor__out,
	output phi_n19__branch_31__ready__0__anchor__out,
	output shl_84__add_85__valid__0__anchor__out,
	output fork_14__icmp_101__ready__0__anchor__out,
	output fork_35__branch_26__data__0__anchor__out,
	output fork_3__branch_21__valid__0__anchor__out,
	output [31 : 0] phi_n11__branch_20__data__0__anchor__out,
	output forkC_45__branchC_47__valid__0__anchor__out,
	output fork_0__load_22__ready__0__anchor__out,
	output fork_35__branch_22__data__0__anchor__out,
	output cst_2__shl_4__valid__0__anchor__out,
	output branchC_52__phiC_34__valid__0__anchor__out,
	output fork_41__branch_43__valid__0__anchor__out,
	output add_59__fork_7__valid__0__anchor__out,
	output fork_35__branch_24__valid__0__anchor__out,
	output fork_9__branch_32__ready__0__anchor__out,
	output [11 : 0] fork_0__add_26__data__0__anchor__out,
	output phiC_33__branchC_52__data__0__anchor__out,
	output forkC_55__branchC_57__valid__0__anchor__out,
	output fork_31__branch_8__ready__0__anchor__out,
	output [5 : 0] branch_7__sink_7__data__0__anchor__out,
	output branch_44__sink_30__valid__0__anchor__out,
	output branch_34__sink_23__valid__0__anchor__out,
	output load_8__MC_A__ready__0__anchor__out,
	output phiC_32__forkC_49__valid__0__anchor__out,
	output branch_21__sink_16__ready__0__anchor__out,
	output branch_40__phi_n23__valid__0__anchor__out,
	output branch_28__Buffer_9__ready__0__anchor__out,
	output fork_31__branch_10__ready__0__anchor__out,
	output branchC_49__phiC_31__ready__0__anchor__out,
	output [5 : 0] branch_18__phi_42__data__0__anchor__out,
	output Buffer_16__phiC_28__data__0__anchor__out,
	output fork_29__branch_2__data__0__anchor__out,
	output cst_24__icmp_101__valid__0__anchor__out,
	output [5 : 0] fork_26__store_3__data__0__anchor__out,
	output w_we1,
	output branch_45__sink_31__ready__0__anchor__out,
	output [31 : 0] branch_20__sink_15__data__0__anchor__out,
	output [31 : 0] branch_40__Buffer_8__data__0__anchor__out,
	output phiC_37__forkC_54__ready__0__anchor__out,
	output [5 : 0] fork_22__branch_24__data__0__anchor__out,
	output alpha__branch_2__valid__0__anchor__out,
	output icmp_96__fork_41__data__0__anchor__out,
	output forkC_49__brCst_block6__ready__0__anchor__out,
	output fork_8__load_66__ready__0__anchor__out,
	output branchC_47__sink_33__data__0__anchor__out,
	output fork_41__branchC_58__valid__0__anchor__out,
	output Buffer_6__phiC_38__ready__0__anchor__out,
	output phi_1__branch_4__valid__0__anchor__out,
	output [31 : 0] branch_38__phi_n27__data__0__anchor__out,
	output fork_34__branchC_51__data__0__anchor__out,
	output forkC_49__branchC_51__data__0__anchor__out,
	output source_15__cst_22__ready__0__anchor__out,
	output phiC_29__phi_3__data__0__anchor__out,
	output source_14__cst_21__data__0__anchor__out,
	output [31 : 0] MC_u2__load_19__data__0__anchor__out,
	output fork_30__branch_5__ready__0__anchor__out,
	output [31 : 0] mul_89__mul_93__data__0__anchor__out,
	output MC_v2__load_22__valid__0__anchor__out,
	output fork_40__branchC_57__data__0__anchor__out,
	output forkC_52__cst_15__ready__0__anchor__out,
	output branch_1__phi_n0__valid__0__anchor__out,
	output [5 : 0] source_3__cst_5__data__0__anchor__out,
	output [31 : 0] mul_23__add_24__data__0__anchor__out,
	output MC_A__load_8__valid__0__anchor__out,
	output source_8__cst_12__valid__0__anchor__out,
	output fork_8__add_73__ready__0__anchor__out,
	output fork_33__branchC_50__valid__0__anchor__out,
	output load_8__add_16__ready__0__anchor__out,
	output [31 : 0] Buffer_5__phi_n7__data__0__anchor__out,
	output [5 : 0] fork_6__icmp_55__data__0__anchor__out,
	output [5 : 0] cst_4__add_29__data__0__anchor__out,
	output Buffer_22__phi_n17__valid__0__anchor__out,
	output fork_1__branch_7__ready__0__anchor__out,
	output [10 : 0] fork_17__shl_25__data__0__anchor__out,
	output load_14__MC_v1__valid__0__anchor__out,
	output fork_38__branch_33__ready__0__anchor__out,
	output fork_30__branch_4__ready__0__anchor__out,
	output branch_37__phi_83__ready__0__anchor__out,
	output [31 : 0] add_94__branch_40__data__0__anchor__out,
	output Buffer_0__phi_77__valid__0__anchor__out,
	output forkC_45__brCst_block2__valid__0__anchor__out,
	output branch_3__sink_3__data__0__anchor__out,
	output Buffer_2__phiC_39__ready__0__anchor__out,
	output MC_x__load_92__ready__0__anchor__out,
	output [31 : 0] branch_1__sink_1__data__0__anchor__out,
	output branchC_54__phiC_36__data__0__anchor__out,
	output [31 : 0] Buffer_8__phi_82__data__0__anchor__out,
	output [5 : 0] fork_3__load_39__data__0__anchor__out,
	output Buffer_26__phi_1__ready__0__anchor__out,
	output branchC_58__phiC_40__ready__0__anchor__out,
	output branch_28__sink_19__ready__0__anchor__out,
	output branch_10__phi_n4__ready__0__anchor__out,
	output branch_32__sink_22__valid__0__anchor__out,
	output [31 : 0] branch_22__Buffer_12__data__0__anchor__out,
	output phi_n9__branch_16__valid__0__anchor__out,
	output fork_42__branch_45__valid__0__anchor__out,
	output branch_29__phi_n19__ready__0__anchor__out,
	output cst_11__add_54__ready__0__anchor__out,
	output branch_25__phi_n14__ready__0__anchor__out,
	output Buffer_1__phi_n0__ready__0__anchor__out,
	output icmp_60__fork_36__ready__0__anchor__out,
	output fork_40__branch_36__ready__0__anchor__out,
	output fork_29__branchC_46__valid__0__anchor__out,
	output phiC_34__forkC_51__data__0__anchor__out,
	output branchC_48__phiC_30__data__0__anchor__out,
	output phi_n8__branch_15__valid__0__anchor__out,
	output branch_19__phi_n17__valid__0__anchor__out,
	output branch_24__Buffer_17__ready__0__anchor__out,
	output fork_40__branch_39__ready__0__anchor__out,
	output Buffer_26__phi_1__valid__0__anchor__out,
	output y_ce0,
	output add_70__store_2__valid__0__anchor__out,
	output cst_22__icmp_96__ready__0__anchor__out,
	output cst_8__branch_14__valid__0__anchor__out,
	output MC_u1__end_0__ready__0__anchor__out,
	output phiC_29__phi_3__ready__0__anchor__out,
	output [31 : 0] u2_dout0,
	output branch_34__sink_23__ready__0__anchor__out,
	output z_we0,
	output [31 : 0] Buffer_1__phi_n0__data__0__anchor__out,
	output branch_11__Buffer_26__ready__0__anchor__out,
	output fork_29__branch_2__valid__0__anchor__out,
	output load_22__MC_v2__ready__0__anchor__out,
	output [31 : 0] phi_n7__branch_10__data__0__anchor__out,
	output branch_33__phi_n21__ready__0__anchor__out,
	output [5 : 0] u2_address0,
	output [5 : 0] branch_45__sink_31__data__0__anchor__out,
	output phi_n16__fork_22__valid__0__anchor__out,
	output branchC_53__Buffer_27__valid__0__anchor__out,
	output icmp_30__fork_31__ready__0__anchor__out,
	output [2 : 0] source_13__cst_20__data__0__anchor__out,
	output fork_17__load_11__valid__0__anchor__out,
	output load_88__MC_A__valid__0__anchor__out,
	output phi_63__fork_8__ready__0__anchor__out,
	output fork_41__branch_41__ready__0__anchor__out,
	output forkC_51__cst_26__valid__0__anchor__out,
	output MC_A__end_0__ready__0__anchor__out,
	output [5 : 0] load_80__MC_w__data__0__anchor__out,
	output [5 : 0] branch_8__phi_n2__data__0__anchor__out,
	output fork_14__icmp_101__valid__0__anchor__out,
	output fork_32__branch_13__valid__0__anchor__out,
	output cst_1__branch_3__ready__0__anchor__out,
	output branch_14__phi_36__ready__0__anchor__out,
	output branch_32__Buffer_10__valid__0__anchor__out,
	output fork_36__branch_27__valid__0__anchor__out,
	output u1_ce1,
	output Buffer_17__phi_n16__ready__0__anchor__out,
	output fork_22__branch_24__valid__0__anchor__out,
	output [5 : 0] fork_2__icmp_33__data__0__anchor__out,
	output branchC_57__phiC_39__valid__0__anchor__out,
	output [5 : 0] source_12__cst_17__data__0__anchor__out,
	output fork_65__phi_83__ready__0__anchor__out,
	output [31 : 0] branch_36__sink_25__data__0__anchor__out,
	output source_1__cst_3__valid__0__anchor__out,
	output cst_12__icmp_55__ready__0__anchor__out,
	output Buffer_11__phi_n22__ready__0__anchor__out,
	output phiC_28__forkC_45__valid__0__anchor__out,
	output branch_33__Buffer_28__valid__0__anchor__out,
	output forkC_52__branchC_54__valid__0__anchor__out,
	output branchC_48__phiC_30__ready__0__anchor__out,
	output fork_29__branch_0__ready__0__anchor__out,
	output [31 : 0] branch_20__phi_n18__data__0__anchor__out,
	output [31 : 0] beta__branch_1__data__0__anchor__out,
	output phi_n23__store_3__ready__0__anchor__out,
	output [31 : 0] load_11__mul_15__data__0__anchor__out,
	output [5 : 0] add_100__fork_14__data__0__anchor__out,
	output Buffer_15__phi_n26__valid__0__anchor__out,
	output load_19__MC_u2__valid__0__anchor__out,
	output fork_65__phi_82__ready__0__anchor__out,
	output fork_34__branch_18__ready__0__anchor__out,
	output [5 : 0] cst_7__icmp_33__data__0__anchor__out,
	output [5 : 0] phi_77__fork_10__data__0__anchor__out,
	output forkC_44__branchC_46__ready__0__anchor__out,
	output fork_27__branch_42__valid__0__anchor__out,
	output add_85__load_88__ready__0__anchor__out,
	output branch_8__phi_n2__ready__0__anchor__out,
	output [31 : 0] phi_n4__branch_13__data__0__anchor__out,
	output [31 : 0] MC_A__load_8__data__0__anchor__out,
	output fork_40__branch_36__data__0__anchor__out,
	output [5 : 0] fork_17__load_11__data__0__anchor__out,
	output branchC_48__Buffer_20__data__0__anchor__out,
	output load_19__MC_u2__ready__0__anchor__out,
	output [31 : 0] branch_31__phi_n20__data__0__anchor__out,
	output alpha_ready_in,
	output phiC_31__forkC_48__data__0__anchor__out,
	output source_16__cst_23__data__0__anchor__out,
	output fork_41__branch_43__data__0__anchor__out,
	output [5 : 0] Buffer_25__phi_3__data__0__anchor__out,
	output beta__branch_1__ready__0__anchor__out,
	output mul_15__add_16__ready__0__anchor__out,
	output fork_36__branch_29__ready__0__anchor__out,
	output [5 : 0] x_address1,
	output source_9__cst_13__data__0__anchor__out,
	output branchC_50__phiC_32__valid__0__anchor__out,
	output branch_12__Buffer_1__ready__0__anchor__out,
	output fork_26__store_3__valid__0__anchor__out,
	output fork_38__branch_32__valid__0__anchor__out,
	output branch_16__sink_11__valid__0__anchor__out,
	output [5 : 0] load_92__MC_x__data__0__anchor__out,
	output fork_35__branchC_52__data__0__anchor__out,
	output branch_0__sink_0__ready__0__anchor__out,
	output branch_0__sink_0__valid__0__anchor__out,
	output phiC_38__phi_77__ready__0__anchor__out,
	output load_69__add_70__valid__0__anchor__out,
	output y_ce1,
	output [31 : 0] branch_10__Buffer_5__data__0__anchor__out,
	output fork_35__branch_25__ready__0__anchor__out,
	output [5 : 0] phi_1__branch_4__data__0__anchor__out,
	output branchC_50__sink_34__data__0__anchor__out,
	output branch_43__phi_n25__ready__0__anchor__out,
	output load_47__mul_48__valid__0__anchor__out,
	output branch_44__sink_30__ready__0__anchor__out,
	output [2 : 0] source_0__cst_2__data__0__anchor__out,
	output [31 : 0] store_3__MC_w__data__0__anchor__out,
	output branch_25__Buffer_22__ready__0__anchor__out,
	output fork_35__branchC_52__ready__0__anchor__out,
	output [31 : 0] cst_25__MC_A__data__0__anchor__out,
	output branchC_57__sink_38__ready__0__anchor__out,
	output phiC_32__phi_36__valid__0__anchor__out,
	output u1_we1,
	output icmp_33__fork_32__ready__0__anchor__out,
	output source_3__cst_5__valid__0__anchor__out,
	output [31 : 0] load_39__branch_17__data__0__anchor__out,
	output Buffer_3__phi_42__valid__0__anchor__out,
	output alpha__branch_2__ready__0__anchor__out,
	output [5 : 0] fork_6__branch_23__data__0__anchor__out,
	output [31 : 0] load_69__add_70__data__0__anchor__out,
	output branch_34__phi_77__ready__0__anchor__out,
	output cst_15__branch_30__ready__0__anchor__out,
	output branchC_50__sink_34__valid__0__anchor__out,
	output branch_42__Buffer_15__ready__0__anchor__out,
	output phi_n10__branch_19__valid__0__anchor__out,
	output forkC_49__cst_9__ready__0__anchor__out,
	output phi_n18__branch_26__valid__0__anchor__out,
	output branch_31__sink_21__valid__0__anchor__out,
	output v1_we0,
	output icmp_30__fork_31__data__0__anchor__out,
	output branch_13__phi_n9__valid__0__anchor__out,
	output [5 : 0] source_5__cst_7__data__0__anchor__out,
	output shl_25__add_26__valid__0__anchor__out,
	output add_32__fork_2__ready__0__anchor__out,
	output phi_n4__branch_13__ready__0__anchor__out,
	output [11 : 0] load_8__MC_A__data__0__anchor__out,
	output [31 : 0] mul_52__add_53__data__0__anchor__out,
	output Buffer_7__phiC_36__ready__0__anchor__out,
	output fork_11__load_92__valid__0__anchor__out,
	output fork_35__branchC_52__valid__0__anchor__out,
	output fork_41__branchC_58__data__0__anchor__out,
	output branch_19__phi_n17__ready__0__anchor__out,
	output Buffer_14__phi_n5__valid__0__anchor__out,
	output v1_ce1,
	output phiC_40__forkC_57__valid__0__anchor__out,
	output fork_4__load_51__valid__0__anchor__out,
	output [5 : 0] phi_n26__fork_27__data__0__anchor__out,
	output fork_38__branchC_55__ready__0__anchor__out,
	output [5 : 0] cst_5__icmp_30__data__0__anchor__out,
	output [31 : 0] v2_dout1,
	output phi_1__branch_4__ready__0__anchor__out,
	output fork_30__branch_4__valid__0__anchor__out,
	output fork_37__branchC_54__ready__0__anchor__out,
	output branchC_52__phiC_34__ready__0__anchor__out,
	output branch_14__phi_36__valid__0__anchor__out,
	output fork_34__branch_19__valid__0__anchor__out,
	output cst_16__add_73__ready__0__anchor__out,
	output MC_A__end_0__valid__0__anchor__out,
	output [5 : 0] branch_11__sink_8__data__0__anchor__out,
	output [31 : 0] load_51__mul_52__data__0__anchor__out,
	output brCst_block12__fork_40__valid__0__anchor__out,
	output phi_n12__store_1__ready__0__anchor__out,
	output [5 : 0] Buffer_10__phi_63__data__0__anchor__out,
	output fork_8__load_66__valid__0__anchor__out,
	output branch_17__phi_41__ready__0__anchor__out,
	output fork_7__icmp_60__ready__0__anchor__out,
	output load_88__mul_89__valid__0__anchor__out,
	output branch_28__sink_19__valid__0__anchor__out,
	output MC_v1__end_0__data__0__anchor__out,
	output fork_23__branch_25__ready__0__anchor__out,
	output fork_32__branch_13__data__0__anchor__out,
	output forkC_57__cst_28__ready__0__anchor__out,
	output [31 : 0] Buffer_11__phi_n22__data__0__anchor__out,
	output fork_13__branch_41__valid__0__anchor__out,
	output branch_3__phi_3__ready__0__anchor__out,
	output phiC_39__branchC_58__data__0__anchor__out,
	output [31 : 0] branch_22__phi_n12__data__0__anchor__out,
	output [5 : 0] branch_24__Buffer_17__data__0__anchor__out,
	output branchC_49__Buffer_16__valid__0__anchor__out,
	output load_92__mul_93__ready__0__anchor__out,
	output MC_u2__end_0__valid__0__anchor__out,
	output cst_13__add_59__valid__0__anchor__out,
	output A_ce0,
	output [5 : 0] Buffer_0__phi_77__data__0__anchor__out,
	output Buffer_20__phiC_29__data__0__anchor__out,
	output fork_33__branch_14__valid__0__anchor__out,
	output MC_x__end_0__ready__0__anchor__out,
	output load_14__mul_15__ready__0__anchor__out,
	output source_0__cst_2__valid__0__anchor__out,
	output source_7__cst_11__ready__0__anchor__out,
	output source_9__cst_13__valid__0__anchor__out,
	output fork_30__branch_6__data__0__anchor__out,
	output fork_30__branch_3__data__0__anchor__out,
	output phiC_28__phi_1__data__0__anchor__out,
	output z_ce1,
	output forkC_54__branchC_56__ready__0__anchor__out,
	output fork_11__add_95__valid__0__anchor__out,
	output [5 : 0] u1_address0,
	output branch_22__phi_n12__valid__0__anchor__out,
	output [31 : 0] MC_u1__load_11__data__0__anchor__out,
	output fork_0__add_26__valid__0__anchor__out,
	output branchC_50__sink_34__ready__0__anchor__out,
	output fork_35__branch_23__ready__0__anchor__out,
	output branch_21__phi_n16__valid__0__anchor__out,
	output branchC_58__Buffer_2__valid__0__anchor__out,
	output branch_24__phi_n13__valid__0__anchor__out,
	output branch_40__Buffer_8__ready__0__anchor__out,
	output phiC_29__forkC_46__ready__0__anchor__out,
	output [5 : 0] phi_n24__fork_26__data__0__anchor__out,
	output MC_A__load_47__ready__0__anchor__out,
	output branch_45__Buffer_0__ready__0__anchor__out,
	output cst_26__MC_x__valid__0__anchor__out,
	output forkC_48__branchC_50__data__0__anchor__out,
	output fork_31__branch_7__ready__0__anchor__out,
	output [31 : 0] add_53__branch_22__data__0__anchor__out,
	output fork_41__branch_42__data__0__anchor__out,
	output cst_10__shl_43__valid__0__anchor__out,
	output fork_40__branch_38__ready__0__anchor__out,
	output phi_n25__branch_44__valid__0__anchor__out,
	output [31 : 0] MC_x__load_39__data__0__anchor__out,
	output MC_u2__end_0__data__0__anchor__out,
	output branch_36__phi_82__valid__0__anchor__out,
	output [31 : 0] y_dout0,
	output fork_6__branch_23__valid__0__anchor__out,
	output phiC_29__phi_3__valid__0__anchor__out,
	output u1_we0,
	output fork_28__branch_43__valid__0__anchor__out,
	output [5 : 0] Buffer_17__phi_n16__data__0__anchor__out,
	output store_0__MC_A__valid__0__anchor__out,
	output branchC_50__phiC_32__data__0__anchor__out,
	output forkC_53__branchC_55__data__0__anchor__out,
	output phi_n19__branch_31__valid__0__anchor__out,
	output phiC_32__phi_36__data__0__anchor__out,
	output u2_ce1,
	output [31 : 0] phi_n15__branch_29__data__0__anchor__out,
	output beta__branch_1__valid__0__anchor__out,
	output MC_u2__load_19__ready__0__anchor__out,
	output cst_7__icmp_33__ready__0__anchor__out,
	output [2 : 0] source_1__cst_3__data__0__anchor__out,
	output load_88__MC_A__ready__0__anchor__out,
	output fork_20__store_1__valid__0__anchor__out,
	output forkC_53__cst_27__data__0__anchor__out,
	output branch_2__sink_2__ready__0__anchor__out,
	output branch_8__phi_n2__valid__0__anchor__out,
	output fork_40__branch_39__data__0__anchor__out,
	output start_ready,
	output u1_ce0,
	output source_3__cst_5__ready__0__anchor__out,
	output icmp_101__fork_42__ready__0__anchor__out,
	output Buffer_5__phi_n7__valid__0__anchor__out,
	output Buffer_6__phiC_38__data__0__anchor__out,
	output fork_7__icmp_60__valid__0__anchor__out,
	output branch_20__phi_n18__valid__0__anchor__out,
	output phi_n24__fork_26__ready__0__anchor__out,
	output cst_23__add_100__ready__0__anchor__out,
	output [5 : 0] add_29__fork_1__data__0__anchor__out,
	output mul_89__mul_93__valid__0__anchor__out,
	output shl_4__add_5__ready__0__anchor__out,
	output phiC_33__branchC_52__ready__0__anchor__out,
	output [31 : 0] Buffer_13__phi_n10__data__0__anchor__out,
	output [31 : 0] Buffer_18__phi_n18__data__0__anchor__out,
	output fork_32__branch_12__valid__0__anchor__out,
	output branch_39__phi_n26__ready__0__anchor__out,
	output forkC_48__brCst_block5__valid__0__anchor__out,
	output [5 : 0] fork_11__load_92__data__0__anchor__out,
	output branchC_53__Buffer_27__data__0__anchor__out,
	output branch_21__sink_16__valid__0__anchor__out,
	output mul_48__mul_52__ready__0__anchor__out,
	output fork_39__branch_35__ready__0__anchor__out,
	output [5 : 0] branch_45__Buffer_0__data__0__anchor__out,
	output branchC_51__phiC_33__valid__0__anchor__out,
	output add_95__fork_13__ready__0__anchor__out,
	output MC_u1__load_11__valid__0__anchor__out,
	output cst_12__icmp_55__valid__0__anchor__out,
	output load_80__branch_36__valid__0__anchor__out,
	output branch_11__sink_8__valid__0__anchor__out,
	output load_22__MC_v2__valid__0__anchor__out,
	output Buffer_16__phiC_28__ready__0__anchor__out,
	output fork_10__branch_39__valid__0__anchor__out,
	output forkC_52__brCst_block9__ready__0__anchor__out,
	output forkC_57__branchC_59__ready__0__anchor__out,
	output [5 : 0] add_59__fork_7__data__0__anchor__out,
	output phi_n26__fork_27__valid__0__anchor__out,
	output [10 : 0] cst_2__shl_4__data__0__anchor__out,
	output load_8__MC_A__valid__0__anchor__out,
	output branch_0__sink_0__data__0__anchor__out,
	output load_92__MC_x__ready__0__anchor__out,
	output fork_39__branch_35__valid__0__anchor__out,
	output phi_n3__branch_12__ready__0__anchor__out,
	output branch_13__phi_n9__ready__0__anchor__out,
	output load_51__MC_y__valid__0__anchor__out,
	output mul_52__add_53__ready__0__anchor__out,
	output [5 : 0] phi_n2__add_32__data__0__anchor__out,
	output branch_38__sink_27__valid__0__anchor__out,
	output forkC_52__brCst_block9__data__0__anchor__out,
	output branchC_55__phiC_37__valid__0__anchor__out,
	output cst_21__add_95__valid__0__anchor__out,
	output [5 : 0] w_address1,
	output branch_18__phi_42__valid__0__anchor__out,
	output Buffer_24__phi_n11__valid__0__anchor__out,
	output fork_22__add_44__ready__0__anchor__out,
	output Buffer_23__phi_n27__ready__0__anchor__out,
	output store_2__MC_x__ready__0__anchor__out,
	output [5 : 0] branch_34__phi_77__data__0__anchor__out,
	output [31 : 0] w_dout1,
	output MC_v1__end_0__valid__0__anchor__out,
	output branchC_59__Buffer_6__data__0__anchor__out,
	output forkC_55__cst_19__data__0__anchor__out,
	output branchC_55__phiC_37__ready__0__anchor__out,
	output [5 : 0] fork_1__branch_7__data__0__anchor__out,
	output MC_v2__end_0__ready__0__anchor__out,
	output [10 : 0] fork_4__shl_43__data__0__anchor__out,
	output cst_14__icmp_60__ready__0__anchor__out,
	output fork_42__branch_44__data__0__anchor__out,
	output fork_4__shl_43__valid__0__anchor__out,
	output phiC_34__forkC_51__ready__0__anchor__out,
	output icmp_74__fork_38__data__0__anchor__out,
	output Buffer_18__phi_n18__valid__0__anchor__out,
	output source_13__cst_20__ready__0__anchor__out,
	output [31 : 0] A_dout1,
	output branch_9__phi_n3__valid__0__anchor__out,
	output fork_33__branch_15__valid__0__anchor__out,
	output forkC_44__branchC_46__valid__0__anchor__out,
	output phi_n5__fork_17__ready__0__anchor__out,
	output [31 : 0] phi_n9__branch_16__data__0__anchor__out,
	output [5 : 0] load_39__MC_x__data__0__anchor__out,
	output phiC_28__phi_1__valid__0__anchor__out,
	output branchC_58__Buffer_2__data__0__anchor__out,
	output [5 : 0] Buffer_26__phi_1__data__0__anchor__out,
	output fork_9__branch_32__valid__0__anchor__out,
	output MC_v2__end_0__data__0__anchor__out,
	output [5 : 0] phi_42__fork_4__data__0__anchor__out,
	output fork_17__branch_8__valid__0__anchor__out,
	output [5 : 0] fork_7__branch_28__data__0__anchor__out,
	output fork_32__branchC_49__ready__0__anchor__out,
	output source_0__cst_2__ready__0__anchor__out,
	output [31 : 0] phi_n17__fork_23__data__0__anchor__out,
	output brCst_block2__fork_30__data__0__anchor__out,
	output [31 : 0] branch_25__Buffer_22__data__0__anchor__out,
	output phi_n20__branch_33__ready__0__anchor__out,
	output Buffer_4__phi_n6__valid__0__anchor__out,
	output icmp_96__fork_41__valid__0__anchor__out,
	output fork_4__add_54__valid__0__anchor__out,
	output fork_3__load_39__ready__0__anchor__out,
	output phi_3__fork_0__valid__0__anchor__out,
	output brCst_block1__fork_29__ready__0__anchor__out,
	output [31 : 0] branch_29__phi_n19__data__0__anchor__out,
	output branchC_55__Buffer_7__valid__0__anchor__out,
	output phiC_41__ret_0__data__0__anchor__out,
	output Buffer_2__phiC_39__valid__0__anchor__out,
	output mul_93__add_94__ready__0__anchor__out,
	output MC_x__end_0__data__0__anchor__out,
	output phi_n12__store_1__valid__0__anchor__out,
	output source_11__cst_16__valid__0__anchor__out,
	output icmp_55__fork_35__data__0__anchor__out,
	output [5 : 0] z_address1,
	output [31 : 0] phi_n18__branch_26__data__0__anchor__out,
	output branch_23__Buffer_3__valid__0__anchor__out,
	output fork_41__branch_40__valid__0__anchor__out,
	output fork_62__phi_41__valid__0__anchor__out,
	output branch_41__sink_29__ready__0__anchor__out,
	output load_22__mul_23__ready__0__anchor__out,
	output [5 : 0] load_19__MC_u2__data__0__anchor__out,
	output phi_n4__branch_13__valid__0__anchor__out,
	output fork_20__store_1__ready__0__anchor__out,
	output fork_34__branch_21__ready__0__anchor__out,
	output branchC_49__phiC_31__data__0__anchor__out,
	output fork_36__branch_28__ready__0__anchor__out,
	output branch_0__phi_1__valid__0__anchor__out,
	output fork_35__branch_24__data__0__anchor__out,
	output [5 : 0] branch_42__phi_n24__data__0__anchor__out,
	output cst_1__branch_3__valid__0__anchor__out,
	output Buffer_24__phi_n11__ready__0__anchor__out,
	output [31 : 0] branch_40__phi_n23__data__0__anchor__out,
	output branchC_47__sink_33__ready__0__anchor__out,
	output branchC_56__phiC_38__data__0__anchor__out,
	output [5 : 0] add_95__fork_13__data__0__anchor__out,
	output branchC_46__phiC_28__data__0__anchor__out,
	output [5 : 0] cst_6__add_32__data__0__anchor__out,
	output forkC_55__cst_19__valid__0__anchor__out,
	output load_39__MC_x__ready__0__anchor__out,
	output [5 : 0] load_14__MC_v1__data__0__anchor__out,
	output phi_n26__fork_27__ready__0__anchor__out,
	output z_ce0,
	output [5 : 0] fork_14__icmp_101__data__0__anchor__out,
	output [31 : 0] phi_n3__branch_12__data__0__anchor__out,
	output branchC_47__phiC_29__data__0__anchor__out,
	output fork_29__branch_0__valid__0__anchor__out,
	output branchC_46__sink_32__valid__0__anchor__out,
	output phiC_32__forkC_49__data__0__anchor__out,
	output [5 : 0] branch_8__Buffer_14__data__0__anchor__out,
	output [31 : 0] branch_13__Buffer_19__data__0__anchor__out,
	output branch_15__sink_10__valid__0__anchor__out,
	output phiC_36__forkC_53__data__0__anchor__out,
	output add_59__fork_7__ready__0__anchor__out,
	output branch_23__sink_17__valid__0__anchor__out,
	output fork_1__branch_7__valid__0__anchor__out,
	output fork_1__icmp_30__ready__0__anchor__out,
	output cst_4__add_29__valid__0__anchor__out,
	output fork_32__branch_12__ready__0__anchor__out,
	output MC_y__load_51__ready__0__anchor__out,
	output branchC_46__phiC_28__ready__0__anchor__out,
	output phiC_39__branchC_58__valid__0__anchor__out,
	output fork_23__mul_48__ready__0__anchor__out,
	output branchC_55__phiC_37__data__0__anchor__out,
	output phiC_37__forkC_54__data__0__anchor__out,
	output [5 : 0] y_address0,
	output [5 : 0] fork_0__load_22__data__0__anchor__out,
	output phiC_34__forkC_51__valid__0__anchor__out,
	output cst_20__shl_84__ready__0__anchor__out,
	output fork_40__branchC_57__valid__0__anchor__out,
	output [31 : 0] u2_dout1,
	output cst_9__branch_18__valid__0__anchor__out,
	output cst_4__add_29__ready__0__anchor__out,
	output fork_17__shl_4__ready__0__anchor__out,
	output source_10__cst_14__valid__0__anchor__out,
	output fork_30__branch_3__ready__0__anchor__out,
	output icmp_60__fork_36__valid__0__anchor__out,
	output icmp_101__fork_42__valid__0__anchor__out,
	output store_0__MC_A__ready__0__anchor__out,
	output forkC_52__cst_15__data__0__anchor__out,
	output phiC_39__fork_65__data__0__anchor__out,
	output MC_A__load_88__valid__0__anchor__out,
	output forkC_57__branchC_59__data__0__anchor__out,
	output fork_40__branch_39__valid__0__anchor__out,
	output forkC_52__branchC_54__data__0__anchor__out,
	output forkC_44__cst_0__ready__0__anchor__out,
	output beta_ready_in,
	output branch_36__phi_82__ready__0__anchor__out,
	output fork_0__add_26__ready__0__anchor__out,
	output fork_31__branchC_48__data__0__anchor__out,
	output fork_41__branch_40__ready__0__anchor__out,
	output brCst_block11__fork_39__data__0__anchor__out,
	output branch_29__Buffer_24__valid__0__anchor__out,
	output phi_41__add_53__valid__0__anchor__out,
	output fork_39__branchC_56__data__0__anchor__out,
	output [5 : 0] branch_7__Buffer_25__data__0__anchor__out,
	output start_0__forkC_44__ready__0__anchor__out,
	output fork_36__branch_27__ready__0__anchor__out,
	output v1_ce0,
	output fork_22__add_44__valid__0__anchor__out,
	output fork_30__branchC_47__valid__0__anchor__out,
	output branch_30__sink_20__ready__0__anchor__out,
	output [5 : 0] branch_41__Buffer_29__data__0__anchor__out,
	output fork_34__branch_21__valid__0__anchor__out,
	output branch_18__sink_13__ready__0__anchor__out,
	output fork_36__branchC_53__ready__0__anchor__out,
	output phi_n24__fork_26__valid__0__anchor__out,
	output brCst_block11__fork_39__ready__0__anchor__out,
	output [31 : 0] phi_n6__branch_9__data__0__anchor__out,
	output brCst_block1__fork_29__valid__0__anchor__out,
	output add_100__fork_14__valid__0__anchor__out,
	output [31 : 0] phiC_38__Buffer_30__data__0__anchor__out,
	output branch_10__Buffer_5__valid__0__anchor__out,
	output phiC_28__forkC_45__ready__0__anchor__out,
	output v2_ce0,
	output fork_0__load_14__valid__0__anchor__out,
	output [31 : 0] load_22__mul_23__data__0__anchor__out,
	output Buffer_10__phi_63__ready__0__anchor__out,
	output add_44__load_47__valid__0__anchor__out,
	output [5 : 0] add_54__fork_6__data__0__anchor__out,
	output [5 : 0] fork_20__add_59__data__0__anchor__out,
	output cst_8__branch_14__data__0__anchor__out,
	output [31 : 0] fork_28__mul_89__data__0__anchor__out,
	output load_47__MC_A__ready__0__anchor__out,
	output branch_32__Buffer_10__ready__0__anchor__out,
	output forkC_49__branchC_51__ready__0__anchor__out,
	output [31 : 0] Buffer_12__phi_41__data__0__anchor__out,
	output branchC_59__phiC_41__valid__0__anchor__out,
	output fork_0__load_14__ready__0__anchor__out,
	output forkC_55__brCst_block12__ready__0__anchor__out,
	output branch_3__phi_3__valid__0__anchor__out,
	output branch_38__sink_27__ready__0__anchor__out,
	output branch_11__sink_8__ready__0__anchor__out,
	output shl_84__add_85__ready__0__anchor__out,
	output branchC_56__sink_37__data__0__anchor__out,
	output cst_11__add_54__valid__0__anchor__out,
	output cst_6__add_32__ready__0__anchor__out,
	output brCst_block5__fork_33__valid__0__anchor__out,
	output [5 : 0] fork_8__load_66__data__0__anchor__out,
	output brCst_block2__fork_30__ready__0__anchor__out,
	output forkC_45__branchC_47__ready__0__anchor__out,
	output brCst_block6__fork_34__data__0__anchor__out,
	output forkC_45__brCst_block2__data__0__anchor__out,
	output end_out,
	output branch_37__phi_83__valid__0__anchor__out,
	output fork_11__add_85__valid__0__anchor__out,
	output fork_42__branchC_59__ready__0__anchor__out,
	output load_11__mul_15__valid__0__anchor__out,
	output MC_w__end_0__data__0__anchor__out,
	output [5 : 0] branch_23__Buffer_3__data__0__anchor__out,
	output phi_n2__add_32__valid__0__anchor__out,
	output [31 : 0] MC_w__load_80__data__0__anchor__out,
	output fork_2__branch_11__valid__0__anchor__out,
	output fork_36__branch_28__valid__0__anchor__out,
	output load_66__MC_x__ready__0__anchor__out,
	output fork_6__icmp_55__ready__0__anchor__out,
	output [31 : 0] w_dout0,
	output [5 : 0] fork_0__add_29__data__0__anchor__out,
	output fork_14__branch_45__valid__0__anchor__out,
	output shl_4__add_5__valid__0__anchor__out,
	output ret_0__end_0__valid__0__anchor__out,
	output forkC_51__cst_26__data__0__anchor__out,
	output branchC_56__phiC_38__valid__0__anchor__out,
	output [11 : 0] add_5__load_8__data__0__anchor__out,
	output [5 : 0] branch_32__sink_22__data__0__anchor__out,
	output cst_28__MC_w__ready__0__anchor__out,
	output [31 : 0] add_24__store_0__data__0__anchor__out,
	output load_66__add_70__ready__0__anchor__out,
	output fork_36__branch_29__valid__0__anchor__out,
	output fork_37__branch_31__valid__0__anchor__out,
	output Buffer_28__phi_n20__ready__0__anchor__out,
	output [31 : 0] z_dout1,
	output source_2__cst_4__ready__0__anchor__out,
	output cst_26__MC_x__ready__0__anchor__out,
	output add_32__fork_2__valid__0__anchor__out,
	output phi_n20__branch_33__valid__0__anchor__out,
	output Buffer_15__phi_n26__ready__0__anchor__out,
	output [5 : 0] fork_13__icmp_96__data__0__anchor__out,
	output branch_22__Buffer_12__valid__0__anchor__out,
	output fork_33__branch_16__ready__0__anchor__out,
	output fork_39__branch_35__data__0__anchor__out,
	output branch_23__sink_17__ready__0__anchor__out,
	output phi_n3__branch_12__valid__0__anchor__out,
	output v2_we1,
	output branch_24__phi_n13__ready__0__anchor__out,
	output phi_n21__branch_35__ready__0__anchor__out,
	output icmp_33__fork_32__data__0__anchor__out,
	output cst_18__branch_34__data__0__anchor__out,
	output fork_9__icmp_74__valid__0__anchor__out,
	output fork_31__branch_9__ready__0__anchor__out,
	output phiC_33__branchC_52__valid__0__anchor__out,
	output brCst_block12__fork_40__data__0__anchor__out,
	output [31 : 0] store_1__MC_x__data__0__anchor__out,
	output cst_21__add_95__ready__0__anchor__out,
	output [31 : 0] phi_n0__branch_5__data__0__anchor__out,
	output fork_0__add_5__valid__0__anchor__out,
	output fork_40__branch_38__data__0__anchor__out,
	output [31 : 0] branch_5__phi_n6__data__0__anchor__out,
	output [31 : 0] branch_15__sink_10__data__0__anchor__out,
	output MC_y__end_0__data__0__anchor__out,
	output branch_26__Buffer_18__valid__0__anchor__out,
	output phi_83__fork_11__valid__0__anchor__out,
	output fork_39__branch_34__ready__0__anchor__out,
	output branch_8__Buffer_14__ready__0__anchor__out,
	output [31 : 0] phi_n21__branch_35__data__0__anchor__out,
	output [31 : 0] fork_23__mul_48__data__0__anchor__out,
	output branch_42__phi_n24__ready__0__anchor__out,
	output cst_0__branch_0__ready__0__anchor__out,
	output branchC_58__Buffer_2__ready__0__anchor__out,
	output branchC_57__sink_38__valid__0__anchor__out,
	output phi_n17__fork_23__ready__0__anchor__out,
	output fork_41__branchC_58__ready__0__anchor__out,
	output fork_36__branchC_53__data__0__anchor__out,
	output [31 : 0] phi_n19__branch_31__data__0__anchor__out,
	output MC_x__end_0__valid__0__anchor__out,
	output forkC_51__cst_26__ready__0__anchor__out,
	output fork_37__branch_30__valid__0__anchor__out,
	output fork_41__branch_41__valid__0__anchor__out,
	output forkC_46__branchC_48__data__0__anchor__out,
	output [11 : 0] A_address0,
	output Buffer_17__phi_n16__valid__0__anchor__out,
	output fork_31__branch_9__valid__0__anchor__out,
	output icmp_74__fork_38__ready__0__anchor__out,
	output branch_39__sink_28__ready__0__anchor__out,
	output [5 : 0] cst_24__icmp_101__data__0__anchor__out,
	output branch_44__Buffer_11__ready__0__anchor__out,
	output branchC_56__sink_37__ready__0__anchor__out,
	output source_17__cst_24__valid__0__anchor__out,
	output w_ce1,
	output fork_30__branchC_47__data__0__anchor__out,
	output phi_82__add_94__ready__0__anchor__out,
	output y_we0,
	output fork_30__branch_4__data__0__anchor__out,
	output [5 : 0] branch_30__phi_63__data__0__anchor__out,
	output store_3__MC_w__valid__0__anchor__out,
	output branch_7__sink_7__ready__0__anchor__out,
	output [5 : 0] branch_23__sink_17__data__0__anchor__out,
	output cst_27__MC_x__valid__0__anchor__out,
	output fork_32__branchC_49__data__0__anchor__out,
	output source_6__cst_10__ready__0__anchor__out,
	output [31 : 0] MC_A__load_88__data__0__anchor__out,
	output [5 : 0] Buffer_9__phi_36__data__0__anchor__out,
	output [31 : 0] load_8__add_16__data__0__anchor__out,
	output fork_35__branch_26__ready__0__anchor__out,
	output Buffer_4__phi_n6__ready__0__anchor__out,
	output branchC_56__phiC_38__ready__0__anchor__out,
	output mul_89__mul_93__ready__0__anchor__out,
	output [31 : 0] fork_28__branch_43__data__0__anchor__out,
	output [31 : 0] load_88__mul_89__data__0__anchor__out,
	output [5 : 0] y_address1,
	output Buffer_12__phi_41__valid__0__anchor__out,
	output branchC_51__sink_35__data__0__anchor__out,
	output [11 : 0] add_26__store_0__data__0__anchor__out,
	output forkC_45__cst_1__valid__0__anchor__out,
	output brCst_block5__fork_33__ready__0__anchor__out,
	output Buffer_19__phi_n1__ready__0__anchor__out,
	output load_11__MC_u1__valid__0__anchor__out,
	output fork_9__icmp_74__ready__0__anchor__out,
	output branch_26__phi_n15__ready__0__anchor__out,
	output source_12__cst_17__valid__0__anchor__out,
	output [31 : 0] MC_v2__load_22__data__0__anchor__out,
	output Buffer_29__phi_83__ready__0__anchor__out,
	output forkC_48__cst_8__data__0__anchor__out,
	output mul_23__add_24__ready__0__anchor__out,
	output fork_37__branch_31__ready__0__anchor__out,
	output fork_38__branch_33__valid__0__anchor__out,
	output branchC_51__sink_35__valid__0__anchor__out,
	output [11 : 0] shl_25__add_26__data__0__anchor__out,
	output branch_6__phi_n7__valid__0__anchor__out,
	output MC_x__load_66__valid__0__anchor__out,
	output [5 : 0] add_73__fork_9__data__0__anchor__out,
	output [10 : 0] fork_17__shl_4__data__0__anchor__out,
	output ret_0__end_0__data__0__anchor__out,
	output phi_n22__branch_38__ready__0__anchor__out,
	output branchC_46__sink_32__data__0__anchor__out,
	output mul_48__mul_52__valid__0__anchor__out,
	output [5 : 0] v2_address1,
	output fork_32__branch_11__data__0__anchor__out,
	output fork_8__load_69__ready__0__anchor__out,
	output add_16__add_24__ready__0__anchor__out,
	output branch_10__Buffer_5__ready__0__anchor__out,
	output load_14__MC_v1__ready__0__anchor__out,
	output phi_42__fork_4__ready__0__anchor__out,
	output [5 : 0] branch_24__phi_n13__data__0__anchor__out,
	output source_11__cst_16__ready__0__anchor__out,
	output v2_we0,
	output [31 : 0] add_70__store_2__data__0__anchor__out,
	output fork_36__branch_27__data__0__anchor__out,
	output cst_19__branch_37__data__0__anchor__out,
	output branch_30__sink_20__valid__0__anchor__out,
	output [5 : 0] fork_8__load_69__data__0__anchor__out,
	output fork_35__branch_25__data__0__anchor__out,
	output add_73__fork_9__valid__0__anchor__out,
	output fork_26__add_100__valid__0__anchor__out,
	output brCst_block1__fork_29__data__0__anchor__out,
	output [31 : 0] add_16__add_24__data__0__anchor__out,
	output [31 : 0] load_19__mul_23__data__0__anchor__out,
	output fork_32__branch_11__valid__0__anchor__out,
	output [5 : 0] load_66__MC_x__data__0__anchor__out,
	output fork_3__branch_21__ready__0__anchor__out,
	output branch_17__sink_12__valid__0__anchor__out,
	output fork_17__load_19__ready__0__anchor__out,
	output cst_18__branch_34__valid__0__anchor__out,
	output cst_18__branch_34__ready__0__anchor__out,
	output add_100__fork_14__ready__0__anchor__out,
	output fork_30__branch_5__valid__0__anchor__out,
	output fork_34__branch_17__data__0__anchor__out,
	output branch_30__phi_63__ready__0__anchor__out,
	output phiC_39__branchC_58__ready__0__anchor__out,
	output fork_32__branch_13__ready__0__anchor__out,
	output branch_7__sink_7__valid__0__anchor__out,
	output cst_5__icmp_30__ready__0__anchor__out,
	output load_88__mul_89__ready__0__anchor__out,
	output forkC_45__cst_1__data__0__anchor__out,
	output fork_20__add_59__valid__0__anchor__out,
	output [5 : 0] w_address0,
	output [5 : 0] v1_address1,
	output [5 : 0] fork_0__load_14__data__0__anchor__out,
	output add_29__fork_1__valid__0__anchor__out,
	output Buffer_3__phi_42__ready__0__anchor__out,
	output fork_0__add_29__valid__0__anchor__out,
	output [5 : 0] fork_4__add_54__data__0__anchor__out,
	output Buffer_6__phiC_38__valid__0__anchor__out,
	output branch_29__phi_n19__valid__0__anchor__out,
	output source_4__cst_6__data__0__anchor__out,
	output branch_10__phi_n4__valid__0__anchor__out,
	output branchC_53__phiC_35__data__0__anchor__out,
	output phiC_41__ret_0__ready__0__anchor__out,
	output branch_45__Buffer_0__valid__0__anchor__out,
	output branch_19__sink_14__valid__0__anchor__out,
	output fork_38__branchC_55__valid__0__anchor__out,
	output branchC_57__phiC_39__ready__0__anchor__out,
	output source_15__cst_22__valid__0__anchor__out,
	output [31 : 0] z_dout0,
	output brCst_block9__fork_37__data__0__anchor__out,
	output [10 : 0] cst_3__shl_25__data__0__anchor__out,
	output branchC_59__phiC_41__ready__0__anchor__out,
	output [31 : 0] phi_n23__store_3__data__0__anchor__out,
	output load_69__MC_z__valid__0__anchor__out,
	output mul_52__add_53__valid__0__anchor__out,
	output phiC_38__phi_77__data__0__anchor__out,
	output load_19__mul_23__valid__0__anchor__out,
	output add_44__load_47__ready__0__anchor__out,
	output end_valid,
	output [5 : 0] fork_9__icmp_74__data__0__anchor__out,
	output cst_19__branch_37__valid__0__anchor__out,
	output forkC_54__cst_18__valid__0__anchor__out,
	output fork_31__branch_9__data__0__anchor__out,
	output Buffer_2__phiC_39__data__0__anchor__out,
	output fork_36__branch_29__data__0__anchor__out,
	output [31 : 0] A_dout0,
	output [5 : 0] load_11__MC_u1__data__0__anchor__out,
	output phi_n13__fork_20__valid__0__anchor__out,
	output branch_4__phi_n5__ready__0__anchor__out,
	output [5 : 0] Buffer_3__phi_42__data__0__anchor__out,
	output forkC_46__branchC_48__valid__0__anchor__out,
	output cst_10__shl_43__ready__0__anchor__out,
	output branch_27__sink_18__valid__0__anchor__out,
	output fork_31__branch_8__valid__0__anchor__out,
	output source_2__cst_4__data__0__anchor__out,
	output branch_1__sink_1__ready__0__anchor__out,
	output [31 : 0] u1_dout1,
	output fork_0__add_29__ready__0__anchor__out,
	output [5 : 0] branch_3__phi_3__data__0__anchor__out,
	output [31 : 0] branch_13__phi_n9__data__0__anchor__out,
	output branch_31__phi_n20__valid__0__anchor__out,
	output [31 : 0] branch_12__Buffer_1__data__0__anchor__out,
	output branch_42__Buffer_15__valid__0__anchor__out,
	output branch_5__sink_5__valid__0__anchor__out,
	output [31 : 0] store_0__MC_A__data__0__anchor__out,
	output fork_31__branchC_48__ready__0__anchor__out,
	output source_7__cst_11__data__0__anchor__out,
	output Buffer_12__phi_41__ready__0__anchor__out,
	output fork_40__branch_37__valid__0__anchor__out,
	output [31 : 0] v1_dout1,
	output [31 : 0] branch_19__phi_n17__data__0__anchor__out,
	output fork_33__branch_16__valid__0__anchor__out,
	output branchC_53__phiC_35__ready__0__anchor__out,
	output fork_23__branch_25__valid__0__anchor__out,
	output MC_u2__end_0__ready__0__anchor__out,
	output branchC_56__sink_37__valid__0__anchor__out,
	output branch_30__phi_63__valid__0__anchor__out,
	output [5 : 0] fork_8__store_2__data__0__anchor__out,
	output MC_x__load_39__ready__0__anchor__out,
	output phiC_32__phi_36__ready__0__anchor__out,
	output fork_2__icmp_33__ready__0__anchor__out,
	output [31 : 0] branch_26__Buffer_18__data__0__anchor__out,
	output [31 : 0] MC_x__load_66__data__0__anchor__out,
	output branch_41__Buffer_29__valid__0__anchor__out,
	output fork_27__shl_84__valid__0__anchor__out,
	output phiC_36__phi_63__ready__0__anchor__out,
	output cst_22__icmp_96__valid__0__anchor__out,
	output branch_20__phi_n18__ready__0__anchor__out,
	output forkC_46__branchC_48__ready__0__anchor__out,
	output add_73__fork_9__ready__0__anchor__out,
	output [5 : 0] phi_n5__fork_17__data__0__anchor__out,
	output [5 : 0] phi_63__fork_8__data__0__anchor__out,
	output forkC_55__branchC_57__ready__0__anchor__out,
	output phi_n14__branch_27__valid__0__anchor__out,
	output load_51__mul_52__valid__0__anchor__out,
	output Buffer_21__phiC_33__data__0__anchor__out,
	output fork_37__branchC_54__valid__0__anchor__out,
	output branchC_55__Buffer_7__data__0__anchor__out,
	output Buffer_21__phiC_33__ready__0__anchor__out,
	output Buffer_21__phiC_33__valid__0__anchor__out,
	output phi_77__fork_10__valid__0__anchor__out,
	output fork_41__branch_40__data__0__anchor__out,
	output branch_27__Buffer_13__valid__0__anchor__out,
	output store_0__MC_A__valid__1__anchor__out,
	output load_11__mul_15__ready__0__anchor__out,
	output Buffer_0__phi_77__ready__0__anchor__out,
	output forkC_44__cst_0__data__0__anchor__out,
	output store_3__MC_w__ready__0__anchor__out,
	output add_29__fork_1__ready__0__anchor__out
);
	wire Buffer_30_clk;
	wire Buffer_30_rst;
	wire [31 : 0] Buffer_30_in1_data;
	wire Buffer_30_in1_ready;
	wire Buffer_30_in1_valid;
	wire [31 : 0] Buffer_30_out1_data;
	wire Buffer_30_out1_ready;
	wire Buffer_30_out1_valid;
	wire alpha_clk;
	wire alpha_rst;
	wire [31 : 0] alpha_in1_data;
	wire alpha_in1_ready;
	wire alpha_in1_valid;
	wire [31 : 0] alpha_out1_data;
	wire alpha_out1_ready;
	wire alpha_out1_valid;
	wire beta_clk;
	wire beta_rst;
	wire [31 : 0] beta_in1_data;
	wire beta_in1_ready;
	wire beta_in1_valid;
	wire [31 : 0] beta_out1_data;
	wire beta_out1_ready;
	wire beta_out1_valid;
	wire brCst_block1_clk;
	wire brCst_block1_rst;
	wire brCst_block1_in1_data;
	wire brCst_block1_in1_ready;
	wire brCst_block1_in1_valid;
	wire brCst_block1_out1_data;
	wire brCst_block1_out1_ready;
	wire brCst_block1_out1_valid;
	wire cst_0_clk;
	wire cst_0_rst;
	wire cst_0_in1_data;
	wire cst_0_in1_ready;
	wire cst_0_in1_valid;
	wire cst_0_out1_data;
	wire cst_0_out1_ready;
	wire cst_0_out1_valid;
	wire phi_1_clk;
	wire phi_1_rst;
	wire phi_1_in1_data;
	wire phi_1_in1_ready;
	wire phi_1_in1_valid;
	wire [5 : 0] phi_1_in2_data;
	wire phi_1_in2_ready;
	wire phi_1_in2_valid;
	wire [5 : 0] phi_1_in3_data;
	wire phi_1_in3_ready;
	wire phi_1_in3_valid;
	wire [5 : 0] phi_1_out1_data;
	wire phi_1_out1_ready;
	wire phi_1_out1_valid;
	wire brCst_block2_clk;
	wire brCst_block2_rst;
	wire brCst_block2_in1_data;
	wire brCst_block2_in1_ready;
	wire brCst_block2_in1_valid;
	wire brCst_block2_out1_data;
	wire brCst_block2_out1_ready;
	wire brCst_block2_out1_valid;
	wire cst_1_clk;
	wire cst_1_rst;
	wire cst_1_in1_data;
	wire cst_1_in1_ready;
	wire cst_1_in1_valid;
	wire cst_1_out1_data;
	wire cst_1_out1_ready;
	wire cst_1_out1_valid;
	wire phi_3_clk;
	wire phi_3_rst;
	wire phi_3_in1_data;
	wire phi_3_in1_ready;
	wire phi_3_in1_valid;
	wire [5 : 0] phi_3_in2_data;
	wire phi_3_in2_ready;
	wire phi_3_in2_valid;
	wire [5 : 0] phi_3_in3_data;
	wire phi_3_in3_ready;
	wire phi_3_in3_valid;
	wire [5 : 0] phi_3_out1_data;
	wire phi_3_out1_ready;
	wire phi_3_out1_valid;
	wire cst_2_clk;
	wire cst_2_rst;
	wire [2 : 0] cst_2_in1_data;
	wire cst_2_in1_ready;
	wire cst_2_in1_valid;
	wire [2 : 0] cst_2_out1_data;
	wire cst_2_out1_ready;
	wire cst_2_out1_valid;
	wire shl_4_clk;
	wire shl_4_rst;
	wire [10 : 0] shl_4_in1_data;
	wire shl_4_in1_ready;
	wire shl_4_in1_valid;
	wire [10 : 0] shl_4_in2_data;
	wire shl_4_in2_ready;
	wire shl_4_in2_valid;
	wire [10 : 0] shl_4_out1_data;
	wire shl_4_out1_ready;
	wire shl_4_out1_valid;
	wire add_5_clk;
	wire add_5_rst;
	wire [11 : 0] add_5_in1_data;
	wire add_5_in1_ready;
	wire add_5_in1_valid;
	wire [11 : 0] add_5_in2_data;
	wire add_5_in2_ready;
	wire add_5_in2_valid;
	wire [11 : 0] add_5_out1_data;
	wire add_5_out1_ready;
	wire add_5_out1_valid;
	wire load_8_clk;
	wire load_8_rst;
	wire [31 : 0] load_8_in1_data;
	wire load_8_in1_ready;
	wire load_8_in1_valid;
	wire [11 : 0] load_8_in2_data;
	wire load_8_in2_ready;
	wire load_8_in2_valid;
	wire [31 : 0] load_8_out1_data;
	wire load_8_out1_ready;
	wire load_8_out1_valid;
	wire [11 : 0] load_8_out2_data;
	wire load_8_out2_ready;
	wire load_8_out2_valid;
	wire load_11_clk;
	wire load_11_rst;
	wire [31 : 0] load_11_in1_data;
	wire load_11_in1_ready;
	wire load_11_in1_valid;
	wire [5 : 0] load_11_in2_data;
	wire load_11_in2_ready;
	wire load_11_in2_valid;
	wire [31 : 0] load_11_out1_data;
	wire load_11_out1_ready;
	wire load_11_out1_valid;
	wire [5 : 0] load_11_out2_data;
	wire load_11_out2_ready;
	wire load_11_out2_valid;
	wire load_14_clk;
	wire load_14_rst;
	wire [31 : 0] load_14_in1_data;
	wire load_14_in1_ready;
	wire load_14_in1_valid;
	wire [5 : 0] load_14_in2_data;
	wire load_14_in2_ready;
	wire load_14_in2_valid;
	wire [31 : 0] load_14_out1_data;
	wire load_14_out1_ready;
	wire load_14_out1_valid;
	wire [5 : 0] load_14_out2_data;
	wire load_14_out2_ready;
	wire load_14_out2_valid;
	wire mul_15_clk;
	wire mul_15_rst;
	wire [15 : 0] mul_15_in1_data;
	wire mul_15_in1_ready;
	wire mul_15_in1_valid;
	wire [15 : 0] mul_15_in2_data;
	wire mul_15_in2_ready;
	wire mul_15_in2_valid;
	wire [31 : 0] mul_15_out1_data;
	wire mul_15_out1_ready;
	wire mul_15_out1_valid;
	wire add_16_clk;
	wire add_16_rst;
	wire [31 : 0] add_16_in1_data;
	wire add_16_in1_ready;
	wire add_16_in1_valid;
	wire [31 : 0] add_16_in2_data;
	wire add_16_in2_ready;
	wire add_16_in2_valid;
	wire [31 : 0] add_16_out1_data;
	wire add_16_out1_ready;
	wire add_16_out1_valid;
	wire load_19_clk;
	wire load_19_rst;
	wire [31 : 0] load_19_in1_data;
	wire load_19_in1_ready;
	wire load_19_in1_valid;
	wire [5 : 0] load_19_in2_data;
	wire load_19_in2_ready;
	wire load_19_in2_valid;
	wire [31 : 0] load_19_out1_data;
	wire load_19_out1_ready;
	wire load_19_out1_valid;
	wire [5 : 0] load_19_out2_data;
	wire load_19_out2_ready;
	wire load_19_out2_valid;
	wire load_22_clk;
	wire load_22_rst;
	wire [31 : 0] load_22_in1_data;
	wire load_22_in1_ready;
	wire load_22_in1_valid;
	wire [5 : 0] load_22_in2_data;
	wire load_22_in2_ready;
	wire load_22_in2_valid;
	wire [31 : 0] load_22_out1_data;
	wire load_22_out1_ready;
	wire load_22_out1_valid;
	wire [5 : 0] load_22_out2_data;
	wire load_22_out2_ready;
	wire load_22_out2_valid;
	wire mul_23_clk;
	wire mul_23_rst;
	wire [15 : 0] mul_23_in1_data;
	wire mul_23_in1_ready;
	wire mul_23_in1_valid;
	wire [15 : 0] mul_23_in2_data;
	wire mul_23_in2_ready;
	wire mul_23_in2_valid;
	wire [31 : 0] mul_23_out1_data;
	wire mul_23_out1_ready;
	wire mul_23_out1_valid;
	wire add_24_clk;
	wire add_24_rst;
	wire [31 : 0] add_24_in1_data;
	wire add_24_in1_ready;
	wire add_24_in1_valid;
	wire [31 : 0] add_24_in2_data;
	wire add_24_in2_ready;
	wire add_24_in2_valid;
	wire [31 : 0] add_24_out1_data;
	wire add_24_out1_ready;
	wire add_24_out1_valid;
	wire cst_3_clk;
	wire cst_3_rst;
	wire [2 : 0] cst_3_in1_data;
	wire cst_3_in1_ready;
	wire cst_3_in1_valid;
	wire [2 : 0] cst_3_out1_data;
	wire cst_3_out1_ready;
	wire cst_3_out1_valid;
	wire shl_25_clk;
	wire shl_25_rst;
	wire [10 : 0] shl_25_in1_data;
	wire shl_25_in1_ready;
	wire shl_25_in1_valid;
	wire [10 : 0] shl_25_in2_data;
	wire shl_25_in2_ready;
	wire shl_25_in2_valid;
	wire [10 : 0] shl_25_out1_data;
	wire shl_25_out1_ready;
	wire shl_25_out1_valid;
	wire add_26_clk;
	wire add_26_rst;
	wire [11 : 0] add_26_in1_data;
	wire add_26_in1_ready;
	wire add_26_in1_valid;
	wire [11 : 0] add_26_in2_data;
	wire add_26_in2_ready;
	wire add_26_in2_valid;
	wire [11 : 0] add_26_out1_data;
	wire add_26_out1_ready;
	wire add_26_out1_valid;
	wire store_0_clk;
	wire store_0_rst;
	wire [31 : 0] store_0_in1_data;
	wire store_0_in1_ready;
	wire store_0_in1_valid;
	wire [11 : 0] store_0_in2_data;
	wire store_0_in2_ready;
	wire store_0_in2_valid;
	wire [31 : 0] store_0_out1_data;
	wire store_0_out1_ready;
	wire store_0_out1_valid;
	wire [11 : 0] store_0_out2_data;
	wire store_0_out2_ready;
	wire store_0_out2_valid;
	wire cst_4_clk;
	wire cst_4_rst;
	wire cst_4_in1_data;
	wire cst_4_in1_ready;
	wire cst_4_in1_valid;
	wire cst_4_out1_data;
	wire cst_4_out1_ready;
	wire cst_4_out1_valid;
	wire add_29_clk;
	wire add_29_rst;
	wire [5 : 0] add_29_in1_data;
	wire add_29_in1_ready;
	wire add_29_in1_valid;
	wire [5 : 0] add_29_in2_data;
	wire add_29_in2_ready;
	wire add_29_in2_valid;
	wire [5 : 0] add_29_out1_data;
	wire add_29_out1_ready;
	wire add_29_out1_valid;
	wire cst_5_clk;
	wire cst_5_rst;
	wire [5 : 0] cst_5_in1_data;
	wire cst_5_in1_ready;
	wire cst_5_in1_valid;
	wire [5 : 0] cst_5_out1_data;
	wire cst_5_out1_ready;
	wire cst_5_out1_valid;
	wire icmp_30_clk;
	wire icmp_30_rst;
	wire [5 : 0] icmp_30_in1_data;
	wire icmp_30_in1_ready;
	wire icmp_30_in1_valid;
	wire [5 : 0] icmp_30_in2_data;
	wire icmp_30_in2_ready;
	wire icmp_30_in2_valid;
	wire icmp_30_out1_data;
	wire icmp_30_out1_ready;
	wire icmp_30_out1_valid;
	wire cst_6_clk;
	wire cst_6_rst;
	wire cst_6_in1_data;
	wire cst_6_in1_ready;
	wire cst_6_in1_valid;
	wire cst_6_out1_data;
	wire cst_6_out1_ready;
	wire cst_6_out1_valid;
	wire add_32_clk;
	wire add_32_rst;
	wire [5 : 0] add_32_in1_data;
	wire add_32_in1_ready;
	wire add_32_in1_valid;
	wire [5 : 0] add_32_in2_data;
	wire add_32_in2_ready;
	wire add_32_in2_valid;
	wire [5 : 0] add_32_out1_data;
	wire add_32_out1_ready;
	wire add_32_out1_valid;
	wire cst_7_clk;
	wire cst_7_rst;
	wire [5 : 0] cst_7_in1_data;
	wire cst_7_in1_ready;
	wire cst_7_in1_valid;
	wire [5 : 0] cst_7_out1_data;
	wire cst_7_out1_ready;
	wire cst_7_out1_valid;
	wire icmp_33_clk;
	wire icmp_33_rst;
	wire [5 : 0] icmp_33_in1_data;
	wire icmp_33_in1_ready;
	wire icmp_33_in1_valid;
	wire [5 : 0] icmp_33_in2_data;
	wire icmp_33_in2_ready;
	wire icmp_33_in2_valid;
	wire icmp_33_out1_data;
	wire icmp_33_out1_ready;
	wire icmp_33_out1_valid;
	wire brCst_block5_clk;
	wire brCst_block5_rst;
	wire brCst_block5_in1_data;
	wire brCst_block5_in1_ready;
	wire brCst_block5_in1_valid;
	wire brCst_block5_out1_data;
	wire brCst_block5_out1_ready;
	wire brCst_block5_out1_valid;
	wire cst_8_clk;
	wire cst_8_rst;
	wire cst_8_in1_data;
	wire cst_8_in1_ready;
	wire cst_8_in1_valid;
	wire cst_8_out1_data;
	wire cst_8_out1_ready;
	wire cst_8_out1_valid;
	wire phi_36_clk;
	wire phi_36_rst;
	wire phi_36_in1_data;
	wire phi_36_in1_ready;
	wire phi_36_in1_valid;
	wire [5 : 0] phi_36_in2_data;
	wire phi_36_in2_ready;
	wire phi_36_in2_valid;
	wire [5 : 0] phi_36_in3_data;
	wire phi_36_in3_ready;
	wire phi_36_in3_valid;
	wire [5 : 0] phi_36_out1_data;
	wire phi_36_out1_ready;
	wire phi_36_out1_valid;
	wire load_39_clk;
	wire load_39_rst;
	wire [31 : 0] load_39_in1_data;
	wire load_39_in1_ready;
	wire load_39_in1_valid;
	wire [5 : 0] load_39_in2_data;
	wire load_39_in2_ready;
	wire load_39_in2_valid;
	wire [31 : 0] load_39_out1_data;
	wire load_39_out1_ready;
	wire load_39_out1_valid;
	wire [5 : 0] load_39_out2_data;
	wire load_39_out2_ready;
	wire load_39_out2_valid;
	wire brCst_block6_clk;
	wire brCst_block6_rst;
	wire brCst_block6_in1_data;
	wire brCst_block6_in1_ready;
	wire brCst_block6_in1_valid;
	wire brCst_block6_out1_data;
	wire brCst_block6_out1_ready;
	wire brCst_block6_out1_valid;
	wire phi_41_clk;
	wire phi_41_rst;
	wire phi_41_in1_data;
	wire phi_41_in1_ready;
	wire phi_41_in1_valid;
	wire [31 : 0] phi_41_in2_data;
	wire phi_41_in2_ready;
	wire phi_41_in2_valid;
	wire [31 : 0] phi_41_in3_data;
	wire phi_41_in3_ready;
	wire phi_41_in3_valid;
	wire [31 : 0] phi_41_out1_data;
	wire phi_41_out1_ready;
	wire phi_41_out1_valid;
	wire cst_9_clk;
	wire cst_9_rst;
	wire cst_9_in1_data;
	wire cst_9_in1_ready;
	wire cst_9_in1_valid;
	wire cst_9_out1_data;
	wire cst_9_out1_ready;
	wire cst_9_out1_valid;
	wire phi_42_clk;
	wire phi_42_rst;
	wire phi_42_in1_data;
	wire phi_42_in1_ready;
	wire phi_42_in1_valid;
	wire [5 : 0] phi_42_in2_data;
	wire phi_42_in2_ready;
	wire phi_42_in2_valid;
	wire [5 : 0] phi_42_in3_data;
	wire phi_42_in3_ready;
	wire phi_42_in3_valid;
	wire [5 : 0] phi_42_out1_data;
	wire phi_42_out1_ready;
	wire phi_42_out1_valid;
	wire cst_10_clk;
	wire cst_10_rst;
	wire [2 : 0] cst_10_in1_data;
	wire cst_10_in1_ready;
	wire cst_10_in1_valid;
	wire [2 : 0] cst_10_out1_data;
	wire cst_10_out1_ready;
	wire cst_10_out1_valid;
	wire shl_43_clk;
	wire shl_43_rst;
	wire [10 : 0] shl_43_in1_data;
	wire shl_43_in1_ready;
	wire shl_43_in1_valid;
	wire [10 : 0] shl_43_in2_data;
	wire shl_43_in2_ready;
	wire shl_43_in2_valid;
	wire [10 : 0] shl_43_out1_data;
	wire shl_43_out1_ready;
	wire shl_43_out1_valid;
	wire add_44_clk;
	wire add_44_rst;
	wire [11 : 0] add_44_in1_data;
	wire add_44_in1_ready;
	wire add_44_in1_valid;
	wire [11 : 0] add_44_in2_data;
	wire add_44_in2_ready;
	wire add_44_in2_valid;
	wire [11 : 0] add_44_out1_data;
	wire add_44_out1_ready;
	wire add_44_out1_valid;
	wire load_47_clk;
	wire load_47_rst;
	wire [31 : 0] load_47_in1_data;
	wire load_47_in1_ready;
	wire load_47_in1_valid;
	wire [11 : 0] load_47_in2_data;
	wire load_47_in2_ready;
	wire load_47_in2_valid;
	wire [31 : 0] load_47_out1_data;
	wire load_47_out1_ready;
	wire load_47_out1_valid;
	wire [11 : 0] load_47_out2_data;
	wire load_47_out2_ready;
	wire load_47_out2_valid;
	wire mul_48_clk;
	wire mul_48_rst;
	wire [15 : 0] mul_48_in1_data;
	wire mul_48_in1_ready;
	wire mul_48_in1_valid;
	wire [15 : 0] mul_48_in2_data;
	wire mul_48_in2_ready;
	wire mul_48_in2_valid;
	wire [31 : 0] mul_48_out1_data;
	wire mul_48_out1_ready;
	wire mul_48_out1_valid;
	wire load_51_clk;
	wire load_51_rst;
	wire [31 : 0] load_51_in1_data;
	wire load_51_in1_ready;
	wire load_51_in1_valid;
	wire [5 : 0] load_51_in2_data;
	wire load_51_in2_ready;
	wire load_51_in2_valid;
	wire [31 : 0] load_51_out1_data;
	wire load_51_out1_ready;
	wire load_51_out1_valid;
	wire [5 : 0] load_51_out2_data;
	wire load_51_out2_ready;
	wire load_51_out2_valid;
	wire mul_52_clk;
	wire mul_52_rst;
	wire [15 : 0] mul_52_in1_data;
	wire mul_52_in1_ready;
	wire mul_52_in1_valid;
	wire [15 : 0] mul_52_in2_data;
	wire mul_52_in2_ready;
	wire mul_52_in2_valid;
	wire [31 : 0] mul_52_out1_data;
	wire mul_52_out1_ready;
	wire mul_52_out1_valid;
	wire add_53_clk;
	wire add_53_rst;
	wire [31 : 0] add_53_in1_data;
	wire add_53_in1_ready;
	wire add_53_in1_valid;
	wire [31 : 0] add_53_in2_data;
	wire add_53_in2_ready;
	wire add_53_in2_valid;
	wire [31 : 0] add_53_out1_data;
	wire add_53_out1_ready;
	wire add_53_out1_valid;
	wire cst_11_clk;
	wire cst_11_rst;
	wire cst_11_in1_data;
	wire cst_11_in1_ready;
	wire cst_11_in1_valid;
	wire cst_11_out1_data;
	wire cst_11_out1_ready;
	wire cst_11_out1_valid;
	wire add_54_clk;
	wire add_54_rst;
	wire [5 : 0] add_54_in1_data;
	wire add_54_in1_ready;
	wire add_54_in1_valid;
	wire [5 : 0] add_54_in2_data;
	wire add_54_in2_ready;
	wire add_54_in2_valid;
	wire [5 : 0] add_54_out1_data;
	wire add_54_out1_ready;
	wire add_54_out1_valid;
	wire cst_12_clk;
	wire cst_12_rst;
	wire [5 : 0] cst_12_in1_data;
	wire cst_12_in1_ready;
	wire cst_12_in1_valid;
	wire [5 : 0] cst_12_out1_data;
	wire cst_12_out1_ready;
	wire cst_12_out1_valid;
	wire icmp_55_clk;
	wire icmp_55_rst;
	wire [5 : 0] icmp_55_in1_data;
	wire icmp_55_in1_ready;
	wire icmp_55_in1_valid;
	wire [5 : 0] icmp_55_in2_data;
	wire icmp_55_in2_ready;
	wire icmp_55_in2_valid;
	wire icmp_55_out1_data;
	wire icmp_55_out1_ready;
	wire icmp_55_out1_valid;
	wire store_1_clk;
	wire store_1_rst;
	wire [31 : 0] store_1_in1_data;
	wire store_1_in1_ready;
	wire store_1_in1_valid;
	wire [5 : 0] store_1_in2_data;
	wire store_1_in2_ready;
	wire store_1_in2_valid;
	wire [31 : 0] store_1_out1_data;
	wire store_1_out1_ready;
	wire store_1_out1_valid;
	wire [5 : 0] store_1_out2_data;
	wire store_1_out2_ready;
	wire store_1_out2_valid;
	wire cst_13_clk;
	wire cst_13_rst;
	wire cst_13_in1_data;
	wire cst_13_in1_ready;
	wire cst_13_in1_valid;
	wire cst_13_out1_data;
	wire cst_13_out1_ready;
	wire cst_13_out1_valid;
	wire add_59_clk;
	wire add_59_rst;
	wire [5 : 0] add_59_in1_data;
	wire add_59_in1_ready;
	wire add_59_in1_valid;
	wire [5 : 0] add_59_in2_data;
	wire add_59_in2_ready;
	wire add_59_in2_valid;
	wire [5 : 0] add_59_out1_data;
	wire add_59_out1_ready;
	wire add_59_out1_valid;
	wire cst_14_clk;
	wire cst_14_rst;
	wire [5 : 0] cst_14_in1_data;
	wire cst_14_in1_ready;
	wire cst_14_in1_valid;
	wire [5 : 0] cst_14_out1_data;
	wire cst_14_out1_ready;
	wire cst_14_out1_valid;
	wire icmp_60_clk;
	wire icmp_60_rst;
	wire [5 : 0] icmp_60_in1_data;
	wire icmp_60_in1_ready;
	wire icmp_60_in1_valid;
	wire [5 : 0] icmp_60_in2_data;
	wire icmp_60_in2_ready;
	wire icmp_60_in2_valid;
	wire icmp_60_out1_data;
	wire icmp_60_out1_ready;
	wire icmp_60_out1_valid;
	wire brCst_block9_clk;
	wire brCst_block9_rst;
	wire brCst_block9_in1_data;
	wire brCst_block9_in1_ready;
	wire brCst_block9_in1_valid;
	wire brCst_block9_out1_data;
	wire brCst_block9_out1_ready;
	wire brCst_block9_out1_valid;
	wire cst_15_clk;
	wire cst_15_rst;
	wire cst_15_in1_data;
	wire cst_15_in1_ready;
	wire cst_15_in1_valid;
	wire cst_15_out1_data;
	wire cst_15_out1_ready;
	wire cst_15_out1_valid;
	wire phi_63_clk;
	wire phi_63_rst;
	wire phi_63_in1_data;
	wire phi_63_in1_ready;
	wire phi_63_in1_valid;
	wire [5 : 0] phi_63_in2_data;
	wire phi_63_in2_ready;
	wire phi_63_in2_valid;
	wire [5 : 0] phi_63_in3_data;
	wire phi_63_in3_ready;
	wire phi_63_in3_valid;
	wire [5 : 0] phi_63_out1_data;
	wire phi_63_out1_ready;
	wire phi_63_out1_valid;
	wire load_66_clk;
	wire load_66_rst;
	wire [31 : 0] load_66_in1_data;
	wire load_66_in1_ready;
	wire load_66_in1_valid;
	wire [5 : 0] load_66_in2_data;
	wire load_66_in2_ready;
	wire load_66_in2_valid;
	wire [31 : 0] load_66_out1_data;
	wire load_66_out1_ready;
	wire load_66_out1_valid;
	wire [5 : 0] load_66_out2_data;
	wire load_66_out2_ready;
	wire load_66_out2_valid;
	wire load_69_clk;
	wire load_69_rst;
	wire [31 : 0] load_69_in1_data;
	wire load_69_in1_ready;
	wire load_69_in1_valid;
	wire [5 : 0] load_69_in2_data;
	wire load_69_in2_ready;
	wire load_69_in2_valid;
	wire [31 : 0] load_69_out1_data;
	wire load_69_out1_ready;
	wire load_69_out1_valid;
	wire [5 : 0] load_69_out2_data;
	wire load_69_out2_ready;
	wire load_69_out2_valid;
	wire add_70_clk;
	wire add_70_rst;
	wire [31 : 0] add_70_in1_data;
	wire add_70_in1_ready;
	wire add_70_in1_valid;
	wire [31 : 0] add_70_in2_data;
	wire add_70_in2_ready;
	wire add_70_in2_valid;
	wire [31 : 0] add_70_out1_data;
	wire add_70_out1_ready;
	wire add_70_out1_valid;
	wire store_2_clk;
	wire store_2_rst;
	wire [31 : 0] store_2_in1_data;
	wire store_2_in1_ready;
	wire store_2_in1_valid;
	wire [5 : 0] store_2_in2_data;
	wire store_2_in2_ready;
	wire store_2_in2_valid;
	wire [31 : 0] store_2_out1_data;
	wire store_2_out1_ready;
	wire store_2_out1_valid;
	wire [5 : 0] store_2_out2_data;
	wire store_2_out2_ready;
	wire store_2_out2_valid;
	wire cst_16_clk;
	wire cst_16_rst;
	wire cst_16_in1_data;
	wire cst_16_in1_ready;
	wire cst_16_in1_valid;
	wire cst_16_out1_data;
	wire cst_16_out1_ready;
	wire cst_16_out1_valid;
	wire add_73_clk;
	wire add_73_rst;
	wire [5 : 0] add_73_in1_data;
	wire add_73_in1_ready;
	wire add_73_in1_valid;
	wire [5 : 0] add_73_in2_data;
	wire add_73_in2_ready;
	wire add_73_in2_valid;
	wire [5 : 0] add_73_out1_data;
	wire add_73_out1_ready;
	wire add_73_out1_valid;
	wire cst_17_clk;
	wire cst_17_rst;
	wire [5 : 0] cst_17_in1_data;
	wire cst_17_in1_ready;
	wire cst_17_in1_valid;
	wire [5 : 0] cst_17_out1_data;
	wire cst_17_out1_ready;
	wire cst_17_out1_valid;
	wire icmp_74_clk;
	wire icmp_74_rst;
	wire [5 : 0] icmp_74_in1_data;
	wire icmp_74_in1_ready;
	wire icmp_74_in1_valid;
	wire [5 : 0] icmp_74_in2_data;
	wire icmp_74_in2_ready;
	wire icmp_74_in2_valid;
	wire icmp_74_out1_data;
	wire icmp_74_out1_ready;
	wire icmp_74_out1_valid;
	wire brCst_block11_clk;
	wire brCst_block11_rst;
	wire brCst_block11_in1_data;
	wire brCst_block11_in1_ready;
	wire brCst_block11_in1_valid;
	wire brCst_block11_out1_data;
	wire brCst_block11_out1_ready;
	wire brCst_block11_out1_valid;
	wire cst_18_clk;
	wire cst_18_rst;
	wire cst_18_in1_data;
	wire cst_18_in1_ready;
	wire cst_18_in1_valid;
	wire cst_18_out1_data;
	wire cst_18_out1_ready;
	wire cst_18_out1_valid;
	wire phi_77_clk;
	wire phi_77_rst;
	wire phi_77_in1_data;
	wire phi_77_in1_ready;
	wire phi_77_in1_valid;
	wire [5 : 0] phi_77_in2_data;
	wire phi_77_in2_ready;
	wire phi_77_in2_valid;
	wire [5 : 0] phi_77_in3_data;
	wire phi_77_in3_ready;
	wire phi_77_in3_valid;
	wire [5 : 0] phi_77_out1_data;
	wire phi_77_out1_ready;
	wire phi_77_out1_valid;
	wire load_80_clk;
	wire load_80_rst;
	wire [31 : 0] load_80_in1_data;
	wire load_80_in1_ready;
	wire load_80_in1_valid;
	wire [5 : 0] load_80_in2_data;
	wire load_80_in2_ready;
	wire load_80_in2_valid;
	wire [31 : 0] load_80_out1_data;
	wire load_80_out1_ready;
	wire load_80_out1_valid;
	wire [5 : 0] load_80_out2_data;
	wire load_80_out2_ready;
	wire load_80_out2_valid;
	wire brCst_block12_clk;
	wire brCst_block12_rst;
	wire brCst_block12_in1_data;
	wire brCst_block12_in1_ready;
	wire brCst_block12_in1_valid;
	wire brCst_block12_out1_data;
	wire brCst_block12_out1_ready;
	wire brCst_block12_out1_valid;
	wire phi_82_clk;
	wire phi_82_rst;
	wire phi_82_in1_data;
	wire phi_82_in1_ready;
	wire phi_82_in1_valid;
	wire [31 : 0] phi_82_in2_data;
	wire phi_82_in2_ready;
	wire phi_82_in2_valid;
	wire [31 : 0] phi_82_in3_data;
	wire phi_82_in3_ready;
	wire phi_82_in3_valid;
	wire [31 : 0] phi_82_out1_data;
	wire phi_82_out1_ready;
	wire phi_82_out1_valid;
	wire cst_19_clk;
	wire cst_19_rst;
	wire cst_19_in1_data;
	wire cst_19_in1_ready;
	wire cst_19_in1_valid;
	wire cst_19_out1_data;
	wire cst_19_out1_ready;
	wire cst_19_out1_valid;
	wire phi_83_clk;
	wire phi_83_rst;
	wire phi_83_in1_data;
	wire phi_83_in1_ready;
	wire phi_83_in1_valid;
	wire [5 : 0] phi_83_in2_data;
	wire phi_83_in2_ready;
	wire phi_83_in2_valid;
	wire [5 : 0] phi_83_in3_data;
	wire phi_83_in3_ready;
	wire phi_83_in3_valid;
	wire [5 : 0] phi_83_out1_data;
	wire phi_83_out1_ready;
	wire phi_83_out1_valid;
	wire cst_20_clk;
	wire cst_20_rst;
	wire [2 : 0] cst_20_in1_data;
	wire cst_20_in1_ready;
	wire cst_20_in1_valid;
	wire [2 : 0] cst_20_out1_data;
	wire cst_20_out1_ready;
	wire cst_20_out1_valid;
	wire shl_84_clk;
	wire shl_84_rst;
	wire [10 : 0] shl_84_in1_data;
	wire shl_84_in1_ready;
	wire shl_84_in1_valid;
	wire [10 : 0] shl_84_in2_data;
	wire shl_84_in2_ready;
	wire shl_84_in2_valid;
	wire [10 : 0] shl_84_out1_data;
	wire shl_84_out1_ready;
	wire shl_84_out1_valid;
	wire add_85_clk;
	wire add_85_rst;
	wire [11 : 0] add_85_in1_data;
	wire add_85_in1_ready;
	wire add_85_in1_valid;
	wire [11 : 0] add_85_in2_data;
	wire add_85_in2_ready;
	wire add_85_in2_valid;
	wire [11 : 0] add_85_out1_data;
	wire add_85_out1_ready;
	wire add_85_out1_valid;
	wire load_88_clk;
	wire load_88_rst;
	wire [31 : 0] load_88_in1_data;
	wire load_88_in1_ready;
	wire load_88_in1_valid;
	wire [11 : 0] load_88_in2_data;
	wire load_88_in2_ready;
	wire load_88_in2_valid;
	wire [31 : 0] load_88_out1_data;
	wire load_88_out1_ready;
	wire load_88_out1_valid;
	wire [11 : 0] load_88_out2_data;
	wire load_88_out2_ready;
	wire load_88_out2_valid;
	wire mul_89_clk;
	wire mul_89_rst;
	wire [15 : 0] mul_89_in1_data;
	wire mul_89_in1_ready;
	wire mul_89_in1_valid;
	wire [15 : 0] mul_89_in2_data;
	wire mul_89_in2_ready;
	wire mul_89_in2_valid;
	wire [31 : 0] mul_89_out1_data;
	wire mul_89_out1_ready;
	wire mul_89_out1_valid;
	wire load_92_clk;
	wire load_92_rst;
	wire [31 : 0] load_92_in1_data;
	wire load_92_in1_ready;
	wire load_92_in1_valid;
	wire [5 : 0] load_92_in2_data;
	wire load_92_in2_ready;
	wire load_92_in2_valid;
	wire [31 : 0] load_92_out1_data;
	wire load_92_out1_ready;
	wire load_92_out1_valid;
	wire [5 : 0] load_92_out2_data;
	wire load_92_out2_ready;
	wire load_92_out2_valid;
	wire mul_93_clk;
	wire mul_93_rst;
	wire [15 : 0] mul_93_in1_data;
	wire mul_93_in1_ready;
	wire mul_93_in1_valid;
	wire [15 : 0] mul_93_in2_data;
	wire mul_93_in2_ready;
	wire mul_93_in2_valid;
	wire [31 : 0] mul_93_out1_data;
	wire mul_93_out1_ready;
	wire mul_93_out1_valid;
	wire add_94_clk;
	wire add_94_rst;
	wire [31 : 0] add_94_in1_data;
	wire add_94_in1_ready;
	wire add_94_in1_valid;
	wire [31 : 0] add_94_in2_data;
	wire add_94_in2_ready;
	wire add_94_in2_valid;
	wire [31 : 0] add_94_out1_data;
	wire add_94_out1_ready;
	wire add_94_out1_valid;
	wire cst_21_clk;
	wire cst_21_rst;
	wire cst_21_in1_data;
	wire cst_21_in1_ready;
	wire cst_21_in1_valid;
	wire cst_21_out1_data;
	wire cst_21_out1_ready;
	wire cst_21_out1_valid;
	wire add_95_clk;
	wire add_95_rst;
	wire [5 : 0] add_95_in1_data;
	wire add_95_in1_ready;
	wire add_95_in1_valid;
	wire [5 : 0] add_95_in2_data;
	wire add_95_in2_ready;
	wire add_95_in2_valid;
	wire [5 : 0] add_95_out1_data;
	wire add_95_out1_ready;
	wire add_95_out1_valid;
	wire cst_22_clk;
	wire cst_22_rst;
	wire [5 : 0] cst_22_in1_data;
	wire cst_22_in1_ready;
	wire cst_22_in1_valid;
	wire [5 : 0] cst_22_out1_data;
	wire cst_22_out1_ready;
	wire cst_22_out1_valid;
	wire icmp_96_clk;
	wire icmp_96_rst;
	wire [5 : 0] icmp_96_in1_data;
	wire icmp_96_in1_ready;
	wire icmp_96_in1_valid;
	wire [5 : 0] icmp_96_in2_data;
	wire icmp_96_in2_ready;
	wire icmp_96_in2_valid;
	wire icmp_96_out1_data;
	wire icmp_96_out1_ready;
	wire icmp_96_out1_valid;
	wire store_3_clk;
	wire store_3_rst;
	wire [31 : 0] store_3_in1_data;
	wire store_3_in1_ready;
	wire store_3_in1_valid;
	wire [5 : 0] store_3_in2_data;
	wire store_3_in2_ready;
	wire store_3_in2_valid;
	wire [31 : 0] store_3_out1_data;
	wire store_3_out1_ready;
	wire store_3_out1_valid;
	wire [5 : 0] store_3_out2_data;
	wire store_3_out2_ready;
	wire store_3_out2_valid;
	wire cst_23_clk;
	wire cst_23_rst;
	wire cst_23_in1_data;
	wire cst_23_in1_ready;
	wire cst_23_in1_valid;
	wire cst_23_out1_data;
	wire cst_23_out1_ready;
	wire cst_23_out1_valid;
	wire add_100_clk;
	wire add_100_rst;
	wire [5 : 0] add_100_in1_data;
	wire add_100_in1_ready;
	wire add_100_in1_valid;
	wire [5 : 0] add_100_in2_data;
	wire add_100_in2_ready;
	wire add_100_in2_valid;
	wire [5 : 0] add_100_out1_data;
	wire add_100_out1_ready;
	wire add_100_out1_valid;
	wire cst_24_clk;
	wire cst_24_rst;
	wire [5 : 0] cst_24_in1_data;
	wire cst_24_in1_ready;
	wire cst_24_in1_valid;
	wire [5 : 0] cst_24_out1_data;
	wire cst_24_out1_ready;
	wire cst_24_out1_valid;
	wire icmp_101_clk;
	wire icmp_101_rst;
	wire [5 : 0] icmp_101_in1_data;
	wire icmp_101_in1_ready;
	wire icmp_101_in1_valid;
	wire [5 : 0] icmp_101_in2_data;
	wire icmp_101_in2_ready;
	wire icmp_101_in2_valid;
	wire icmp_101_out1_data;
	wire icmp_101_out1_ready;
	wire icmp_101_out1_valid;
	wire ret_0_clk;
	wire ret_0_rst;
	wire ret_0_in1_data;
	wire ret_0_in1_ready;
	wire ret_0_in1_valid;
	wire ret_0_out1_data;
	wire ret_0_out1_ready;
	wire ret_0_out1_valid;
	wire phi_n0_clk;
	wire phi_n0_rst;
	wire [31 : 0] phi_n0_in1_data;
	wire phi_n0_in1_ready;
	wire phi_n0_in1_valid;
	wire [31 : 0] phi_n0_in2_data;
	wire phi_n0_in2_ready;
	wire phi_n0_in2_valid;
	wire [31 : 0] phi_n0_out1_data;
	wire phi_n0_out1_ready;
	wire phi_n0_out1_valid;
	wire phi_n1_clk;
	wire phi_n1_rst;
	wire [31 : 0] phi_n1_in1_data;
	wire phi_n1_in1_ready;
	wire phi_n1_in1_valid;
	wire [31 : 0] phi_n1_in2_data;
	wire phi_n1_in2_ready;
	wire phi_n1_in2_valid;
	wire [31 : 0] phi_n1_out1_data;
	wire phi_n1_out1_ready;
	wire phi_n1_out1_valid;
	wire phi_n2_clk;
	wire phi_n2_rst;
	wire [5 : 0] phi_n2_in1_data;
	wire phi_n2_in1_ready;
	wire phi_n2_in1_valid;
	wire [5 : 0] phi_n2_out1_data;
	wire phi_n2_out1_ready;
	wire phi_n2_out1_valid;
	wire phi_n3_clk;
	wire phi_n3_rst;
	wire [31 : 0] phi_n3_in1_data;
	wire phi_n3_in1_ready;
	wire phi_n3_in1_valid;
	wire [31 : 0] phi_n3_out1_data;
	wire phi_n3_out1_ready;
	wire phi_n3_out1_valid;
	wire phi_n4_clk;
	wire phi_n4_rst;
	wire [31 : 0] phi_n4_in1_data;
	wire phi_n4_in1_ready;
	wire phi_n4_in1_valid;
	wire [31 : 0] phi_n4_out1_data;
	wire phi_n4_out1_ready;
	wire phi_n4_out1_valid;
	wire phi_n5_clk;
	wire phi_n5_rst;
	wire [5 : 0] phi_n5_in1_data;
	wire phi_n5_in1_ready;
	wire phi_n5_in1_valid;
	wire [5 : 0] phi_n5_in2_data;
	wire phi_n5_in2_ready;
	wire phi_n5_in2_valid;
	wire [5 : 0] phi_n5_out1_data;
	wire phi_n5_out1_ready;
	wire phi_n5_out1_valid;
	wire phi_n6_clk;
	wire phi_n6_rst;
	wire [31 : 0] phi_n6_in1_data;
	wire phi_n6_in1_ready;
	wire phi_n6_in1_valid;
	wire [31 : 0] phi_n6_in2_data;
	wire phi_n6_in2_ready;
	wire phi_n6_in2_valid;
	wire [31 : 0] phi_n6_out1_data;
	wire phi_n6_out1_ready;
	wire phi_n6_out1_valid;
	wire phi_n7_clk;
	wire phi_n7_rst;
	wire [31 : 0] phi_n7_in1_data;
	wire phi_n7_in1_ready;
	wire phi_n7_in1_valid;
	wire [31 : 0] phi_n7_in2_data;
	wire phi_n7_in2_ready;
	wire phi_n7_in2_valid;
	wire [31 : 0] phi_n7_out1_data;
	wire phi_n7_out1_ready;
	wire phi_n7_out1_valid;
	wire phi_n8_clk;
	wire phi_n8_rst;
	wire [31 : 0] phi_n8_in1_data;
	wire phi_n8_in1_ready;
	wire phi_n8_in1_valid;
	wire [31 : 0] phi_n8_out1_data;
	wire phi_n8_out1_ready;
	wire phi_n8_out1_valid;
	wire phi_n9_clk;
	wire phi_n9_rst;
	wire [31 : 0] phi_n9_in1_data;
	wire phi_n9_in1_ready;
	wire phi_n9_in1_valid;
	wire [31 : 0] phi_n9_out1_data;
	wire phi_n9_out1_ready;
	wire phi_n9_out1_valid;
	wire phi_n10_clk;
	wire phi_n10_rst;
	wire [31 : 0] phi_n10_in1_data;
	wire phi_n10_in1_ready;
	wire phi_n10_in1_valid;
	wire [31 : 0] phi_n10_in2_data;
	wire phi_n10_in2_ready;
	wire phi_n10_in2_valid;
	wire [31 : 0] phi_n10_out1_data;
	wire phi_n10_out1_ready;
	wire phi_n10_out1_valid;
	wire phi_n11_clk;
	wire phi_n11_rst;
	wire [31 : 0] phi_n11_in1_data;
	wire phi_n11_in1_ready;
	wire phi_n11_in1_valid;
	wire [31 : 0] phi_n11_in2_data;
	wire phi_n11_in2_ready;
	wire phi_n11_in2_valid;
	wire [31 : 0] phi_n11_out1_data;
	wire phi_n11_out1_ready;
	wire phi_n11_out1_valid;
	wire phi_n12_clk;
	wire phi_n12_rst;
	wire [31 : 0] phi_n12_in1_data;
	wire phi_n12_in1_ready;
	wire phi_n12_in1_valid;
	wire [31 : 0] phi_n12_out1_data;
	wire phi_n12_out1_ready;
	wire phi_n12_out1_valid;
	wire phi_n13_clk;
	wire phi_n13_rst;
	wire [5 : 0] phi_n13_in1_data;
	wire phi_n13_in1_ready;
	wire phi_n13_in1_valid;
	wire [5 : 0] phi_n13_out1_data;
	wire phi_n13_out1_ready;
	wire phi_n13_out1_valid;
	wire phi_n14_clk;
	wire phi_n14_rst;
	wire [31 : 0] phi_n14_in1_data;
	wire phi_n14_in1_ready;
	wire phi_n14_in1_valid;
	wire [31 : 0] phi_n14_out1_data;
	wire phi_n14_out1_ready;
	wire phi_n14_out1_valid;
	wire phi_n15_clk;
	wire phi_n15_rst;
	wire [31 : 0] phi_n15_in1_data;
	wire phi_n15_in1_ready;
	wire phi_n15_in1_valid;
	wire [31 : 0] phi_n15_out1_data;
	wire phi_n15_out1_ready;
	wire phi_n15_out1_valid;
	wire phi_n16_clk;
	wire phi_n16_rst;
	wire [5 : 0] phi_n16_in1_data;
	wire phi_n16_in1_ready;
	wire phi_n16_in1_valid;
	wire [5 : 0] phi_n16_in2_data;
	wire phi_n16_in2_ready;
	wire phi_n16_in2_valid;
	wire [5 : 0] phi_n16_out1_data;
	wire phi_n16_out1_ready;
	wire phi_n16_out1_valid;
	wire phi_n17_clk;
	wire phi_n17_rst;
	wire [31 : 0] phi_n17_in1_data;
	wire phi_n17_in1_ready;
	wire phi_n17_in1_valid;
	wire [31 : 0] phi_n17_in2_data;
	wire phi_n17_in2_ready;
	wire phi_n17_in2_valid;
	wire [31 : 0] phi_n17_out1_data;
	wire phi_n17_out1_ready;
	wire phi_n17_out1_valid;
	wire phi_n18_clk;
	wire phi_n18_rst;
	wire [31 : 0] phi_n18_in1_data;
	wire phi_n18_in1_ready;
	wire phi_n18_in1_valid;
	wire [31 : 0] phi_n18_in2_data;
	wire phi_n18_in2_ready;
	wire phi_n18_in2_valid;
	wire [31 : 0] phi_n18_out1_data;
	wire phi_n18_out1_ready;
	wire phi_n18_out1_valid;
	wire phi_n19_clk;
	wire phi_n19_rst;
	wire [31 : 0] phi_n19_in1_data;
	wire phi_n19_in1_ready;
	wire phi_n19_in1_valid;
	wire [31 : 0] phi_n19_out1_data;
	wire phi_n19_out1_ready;
	wire phi_n19_out1_valid;
	wire phi_n20_clk;
	wire phi_n20_rst;
	wire [31 : 0] phi_n20_in1_data;
	wire phi_n20_in1_ready;
	wire phi_n20_in1_valid;
	wire [31 : 0] phi_n20_in2_data;
	wire phi_n20_in2_ready;
	wire phi_n20_in2_valid;
	wire [31 : 0] phi_n20_out1_data;
	wire phi_n20_out1_ready;
	wire phi_n20_out1_valid;
	wire phi_n21_clk;
	wire phi_n21_rst;
	wire [31 : 0] phi_n21_in1_data;
	wire phi_n21_in1_ready;
	wire phi_n21_in1_valid;
	wire [31 : 0] phi_n21_out1_data;
	wire phi_n21_out1_ready;
	wire phi_n21_out1_valid;
	wire phi_n22_clk;
	wire phi_n22_rst;
	wire [31 : 0] phi_n22_in1_data;
	wire phi_n22_in1_ready;
	wire phi_n22_in1_valid;
	wire [31 : 0] phi_n22_in2_data;
	wire phi_n22_in2_ready;
	wire phi_n22_in2_valid;
	wire [31 : 0] phi_n22_out1_data;
	wire phi_n22_out1_ready;
	wire phi_n22_out1_valid;
	wire phi_n23_clk;
	wire phi_n23_rst;
	wire [31 : 0] phi_n23_in1_data;
	wire phi_n23_in1_ready;
	wire phi_n23_in1_valid;
	wire [31 : 0] phi_n23_out1_data;
	wire phi_n23_out1_ready;
	wire phi_n23_out1_valid;
	wire phi_n24_clk;
	wire phi_n24_rst;
	wire [5 : 0] phi_n24_in1_data;
	wire phi_n24_in1_ready;
	wire phi_n24_in1_valid;
	wire [5 : 0] phi_n24_out1_data;
	wire phi_n24_out1_ready;
	wire phi_n24_out1_valid;
	wire phi_n25_clk;
	wire phi_n25_rst;
	wire [31 : 0] phi_n25_in1_data;
	wire phi_n25_in1_ready;
	wire phi_n25_in1_valid;
	wire [31 : 0] phi_n25_out1_data;
	wire phi_n25_out1_ready;
	wire phi_n25_out1_valid;
	wire phi_n26_clk;
	wire phi_n26_rst;
	wire [5 : 0] phi_n26_in1_data;
	wire phi_n26_in1_ready;
	wire phi_n26_in1_valid;
	wire [5 : 0] phi_n26_in2_data;
	wire phi_n26_in2_ready;
	wire phi_n26_in2_valid;
	wire [5 : 0] phi_n26_out1_data;
	wire phi_n26_out1_ready;
	wire phi_n26_out1_valid;
	wire phi_n27_clk;
	wire phi_n27_rst;
	wire [31 : 0] phi_n27_in1_data;
	wire phi_n27_in1_ready;
	wire phi_n27_in1_valid;
	wire [31 : 0] phi_n27_in2_data;
	wire phi_n27_in2_ready;
	wire phi_n27_in2_valid;
	wire [31 : 0] phi_n27_out1_data;
	wire phi_n27_out1_ready;
	wire phi_n27_out1_valid;
	wire fork_0_clk;
	wire fork_0_rst;
	wire [5 : 0] fork_0_in1_data;
	wire fork_0_in1_ready;
	wire fork_0_in1_valid;
	wire [5 : 0] fork_0_out1_data;
	wire fork_0_out1_ready;
	wire fork_0_out1_valid;
	wire [5 : 0] fork_0_out2_data;
	wire fork_0_out2_ready;
	wire fork_0_out2_valid;
	wire [5 : 0] fork_0_out3_data;
	wire fork_0_out3_ready;
	wire fork_0_out3_valid;
	wire [5 : 0] fork_0_out4_data;
	wire fork_0_out4_ready;
	wire fork_0_out4_valid;
	wire [5 : 0] fork_0_out5_data;
	wire fork_0_out5_ready;
	wire fork_0_out5_valid;
	wire fork_1_clk;
	wire fork_1_rst;
	wire [5 : 0] fork_1_in1_data;
	wire fork_1_in1_ready;
	wire fork_1_in1_valid;
	wire [5 : 0] fork_1_out1_data;
	wire fork_1_out1_ready;
	wire fork_1_out1_valid;
	wire [5 : 0] fork_1_out2_data;
	wire fork_1_out2_ready;
	wire fork_1_out2_valid;
	wire fork_2_clk;
	wire fork_2_rst;
	wire [5 : 0] fork_2_in1_data;
	wire fork_2_in1_ready;
	wire fork_2_in1_valid;
	wire [5 : 0] fork_2_out1_data;
	wire fork_2_out1_ready;
	wire fork_2_out1_valid;
	wire [5 : 0] fork_2_out2_data;
	wire fork_2_out2_ready;
	wire fork_2_out2_valid;
	wire fork_3_clk;
	wire fork_3_rst;
	wire [5 : 0] fork_3_in1_data;
	wire fork_3_in1_ready;
	wire fork_3_in1_valid;
	wire [5 : 0] fork_3_out1_data;
	wire fork_3_out1_ready;
	wire fork_3_out1_valid;
	wire [5 : 0] fork_3_out2_data;
	wire fork_3_out2_ready;
	wire fork_3_out2_valid;
	wire fork_4_clk;
	wire fork_4_rst;
	wire [5 : 0] fork_4_in1_data;
	wire fork_4_in1_ready;
	wire fork_4_in1_valid;
	wire [5 : 0] fork_4_out1_data;
	wire fork_4_out1_ready;
	wire fork_4_out1_valid;
	wire [5 : 0] fork_4_out2_data;
	wire fork_4_out2_ready;
	wire fork_4_out2_valid;
	wire [5 : 0] fork_4_out3_data;
	wire fork_4_out3_ready;
	wire fork_4_out3_valid;
	wire fork_6_clk;
	wire fork_6_rst;
	wire [5 : 0] fork_6_in1_data;
	wire fork_6_in1_ready;
	wire fork_6_in1_valid;
	wire [5 : 0] fork_6_out1_data;
	wire fork_6_out1_ready;
	wire fork_6_out1_valid;
	wire [5 : 0] fork_6_out2_data;
	wire fork_6_out2_ready;
	wire fork_6_out2_valid;
	wire fork_7_clk;
	wire fork_7_rst;
	wire [5 : 0] fork_7_in1_data;
	wire fork_7_in1_ready;
	wire fork_7_in1_valid;
	wire [5 : 0] fork_7_out1_data;
	wire fork_7_out1_ready;
	wire fork_7_out1_valid;
	wire [5 : 0] fork_7_out2_data;
	wire fork_7_out2_ready;
	wire fork_7_out2_valid;
	wire fork_8_clk;
	wire fork_8_rst;
	wire [5 : 0] fork_8_in1_data;
	wire fork_8_in1_ready;
	wire fork_8_in1_valid;
	wire [5 : 0] fork_8_out1_data;
	wire fork_8_out1_ready;
	wire fork_8_out1_valid;
	wire [5 : 0] fork_8_out2_data;
	wire fork_8_out2_ready;
	wire fork_8_out2_valid;
	wire [5 : 0] fork_8_out3_data;
	wire fork_8_out3_ready;
	wire fork_8_out3_valid;
	wire [5 : 0] fork_8_out4_data;
	wire fork_8_out4_ready;
	wire fork_8_out4_valid;
	wire fork_9_clk;
	wire fork_9_rst;
	wire [5 : 0] fork_9_in1_data;
	wire fork_9_in1_ready;
	wire fork_9_in1_valid;
	wire [5 : 0] fork_9_out1_data;
	wire fork_9_out1_ready;
	wire fork_9_out1_valid;
	wire [5 : 0] fork_9_out2_data;
	wire fork_9_out2_ready;
	wire fork_9_out2_valid;
	wire fork_10_clk;
	wire fork_10_rst;
	wire [5 : 0] fork_10_in1_data;
	wire fork_10_in1_ready;
	wire fork_10_in1_valid;
	wire [5 : 0] fork_10_out1_data;
	wire fork_10_out1_ready;
	wire fork_10_out1_valid;
	wire [5 : 0] fork_10_out2_data;
	wire fork_10_out2_ready;
	wire fork_10_out2_valid;
	wire fork_11_clk;
	wire fork_11_rst;
	wire [5 : 0] fork_11_in1_data;
	wire fork_11_in1_ready;
	wire fork_11_in1_valid;
	wire [5 : 0] fork_11_out1_data;
	wire fork_11_out1_ready;
	wire fork_11_out1_valid;
	wire [5 : 0] fork_11_out2_data;
	wire fork_11_out2_ready;
	wire fork_11_out2_valid;
	wire [5 : 0] fork_11_out3_data;
	wire fork_11_out3_ready;
	wire fork_11_out3_valid;
	wire fork_13_clk;
	wire fork_13_rst;
	wire [5 : 0] fork_13_in1_data;
	wire fork_13_in1_ready;
	wire fork_13_in1_valid;
	wire [5 : 0] fork_13_out1_data;
	wire fork_13_out1_ready;
	wire fork_13_out1_valid;
	wire [5 : 0] fork_13_out2_data;
	wire fork_13_out2_ready;
	wire fork_13_out2_valid;
	wire fork_14_clk;
	wire fork_14_rst;
	wire [5 : 0] fork_14_in1_data;
	wire fork_14_in1_ready;
	wire fork_14_in1_valid;
	wire [5 : 0] fork_14_out1_data;
	wire fork_14_out1_ready;
	wire fork_14_out1_valid;
	wire [5 : 0] fork_14_out2_data;
	wire fork_14_out2_ready;
	wire fork_14_out2_valid;
	wire fork_17_clk;
	wire fork_17_rst;
	wire [5 : 0] fork_17_in1_data;
	wire fork_17_in1_ready;
	wire fork_17_in1_valid;
	wire [5 : 0] fork_17_out1_data;
	wire fork_17_out1_ready;
	wire fork_17_out1_valid;
	wire [5 : 0] fork_17_out2_data;
	wire fork_17_out2_ready;
	wire fork_17_out2_valid;
	wire [5 : 0] fork_17_out3_data;
	wire fork_17_out3_ready;
	wire fork_17_out3_valid;
	wire [5 : 0] fork_17_out4_data;
	wire fork_17_out4_ready;
	wire fork_17_out4_valid;
	wire [5 : 0] fork_17_out5_data;
	wire fork_17_out5_ready;
	wire fork_17_out5_valid;
	wire fork_20_clk;
	wire fork_20_rst;
	wire [5 : 0] fork_20_in1_data;
	wire fork_20_in1_ready;
	wire fork_20_in1_valid;
	wire [5 : 0] fork_20_out1_data;
	wire fork_20_out1_ready;
	wire fork_20_out1_valid;
	wire [5 : 0] fork_20_out2_data;
	wire fork_20_out2_ready;
	wire fork_20_out2_valid;
	wire fork_22_clk;
	wire fork_22_rst;
	wire [5 : 0] fork_22_in1_data;
	wire fork_22_in1_ready;
	wire fork_22_in1_valid;
	wire [5 : 0] fork_22_out1_data;
	wire fork_22_out1_ready;
	wire fork_22_out1_valid;
	wire [5 : 0] fork_22_out2_data;
	wire fork_22_out2_ready;
	wire fork_22_out2_valid;
	wire fork_23_clk;
	wire fork_23_rst;
	wire [31 : 0] fork_23_in1_data;
	wire fork_23_in1_ready;
	wire fork_23_in1_valid;
	wire [31 : 0] fork_23_out1_data;
	wire fork_23_out1_ready;
	wire fork_23_out1_valid;
	wire [31 : 0] fork_23_out2_data;
	wire fork_23_out2_ready;
	wire fork_23_out2_valid;
	wire fork_26_clk;
	wire fork_26_rst;
	wire [5 : 0] fork_26_in1_data;
	wire fork_26_in1_ready;
	wire fork_26_in1_valid;
	wire [5 : 0] fork_26_out1_data;
	wire fork_26_out1_ready;
	wire fork_26_out1_valid;
	wire [5 : 0] fork_26_out2_data;
	wire fork_26_out2_ready;
	wire fork_26_out2_valid;
	wire fork_27_clk;
	wire fork_27_rst;
	wire [5 : 0] fork_27_in1_data;
	wire fork_27_in1_ready;
	wire fork_27_in1_valid;
	wire [5 : 0] fork_27_out1_data;
	wire fork_27_out1_ready;
	wire fork_27_out1_valid;
	wire [5 : 0] fork_27_out2_data;
	wire fork_27_out2_ready;
	wire fork_27_out2_valid;
	wire fork_28_clk;
	wire fork_28_rst;
	wire [31 : 0] fork_28_in1_data;
	wire fork_28_in1_ready;
	wire fork_28_in1_valid;
	wire [31 : 0] fork_28_out1_data;
	wire fork_28_out1_ready;
	wire fork_28_out1_valid;
	wire [31 : 0] fork_28_out2_data;
	wire fork_28_out2_ready;
	wire fork_28_out2_valid;
	wire branch_0_clk;
	wire branch_0_rst;
	wire branch_0_in1_data;
	wire branch_0_in1_ready;
	wire branch_0_in1_valid;
	wire branch_0_in2_data;
	wire branch_0_in2_ready;
	wire branch_0_in2_valid;
	wire branch_0_out1_data;
	wire branch_0_out1_ready;
	wire branch_0_out1_valid;
	wire branch_0_out2_data;
	wire branch_0_out2_ready;
	wire branch_0_out2_valid;
	wire branch_1_clk;
	wire branch_1_rst;
	wire [31 : 0] branch_1_in1_data;
	wire branch_1_in1_ready;
	wire branch_1_in1_valid;
	wire branch_1_in2_data;
	wire branch_1_in2_ready;
	wire branch_1_in2_valid;
	wire [31 : 0] branch_1_out1_data;
	wire branch_1_out1_ready;
	wire branch_1_out1_valid;
	wire [31 : 0] branch_1_out2_data;
	wire branch_1_out2_ready;
	wire branch_1_out2_valid;
	wire branch_2_clk;
	wire branch_2_rst;
	wire [31 : 0] branch_2_in1_data;
	wire branch_2_in1_ready;
	wire branch_2_in1_valid;
	wire branch_2_in2_data;
	wire branch_2_in2_ready;
	wire branch_2_in2_valid;
	wire [31 : 0] branch_2_out1_data;
	wire branch_2_out1_ready;
	wire branch_2_out1_valid;
	wire [31 : 0] branch_2_out2_data;
	wire branch_2_out2_ready;
	wire branch_2_out2_valid;
	wire fork_29_clk;
	wire fork_29_rst;
	wire fork_29_in1_data;
	wire fork_29_in1_ready;
	wire fork_29_in1_valid;
	wire fork_29_out1_data;
	wire fork_29_out1_ready;
	wire fork_29_out1_valid;
	wire fork_29_out2_data;
	wire fork_29_out2_ready;
	wire fork_29_out2_valid;
	wire fork_29_out3_data;
	wire fork_29_out3_ready;
	wire fork_29_out3_valid;
	wire fork_29_out4_data;
	wire fork_29_out4_ready;
	wire fork_29_out4_valid;
	wire branch_3_clk;
	wire branch_3_rst;
	wire branch_3_in1_data;
	wire branch_3_in1_ready;
	wire branch_3_in1_valid;
	wire branch_3_in2_data;
	wire branch_3_in2_ready;
	wire branch_3_in2_valid;
	wire branch_3_out1_data;
	wire branch_3_out1_ready;
	wire branch_3_out1_valid;
	wire branch_3_out2_data;
	wire branch_3_out2_ready;
	wire branch_3_out2_valid;
	wire branch_4_clk;
	wire branch_4_rst;
	wire [5 : 0] branch_4_in1_data;
	wire branch_4_in1_ready;
	wire branch_4_in1_valid;
	wire branch_4_in2_data;
	wire branch_4_in2_ready;
	wire branch_4_in2_valid;
	wire [5 : 0] branch_4_out1_data;
	wire branch_4_out1_ready;
	wire branch_4_out1_valid;
	wire [5 : 0] branch_4_out2_data;
	wire branch_4_out2_ready;
	wire branch_4_out2_valid;
	wire branch_5_clk;
	wire branch_5_rst;
	wire [31 : 0] branch_5_in1_data;
	wire branch_5_in1_ready;
	wire branch_5_in1_valid;
	wire branch_5_in2_data;
	wire branch_5_in2_ready;
	wire branch_5_in2_valid;
	wire [31 : 0] branch_5_out1_data;
	wire branch_5_out1_ready;
	wire branch_5_out1_valid;
	wire [31 : 0] branch_5_out2_data;
	wire branch_5_out2_ready;
	wire branch_5_out2_valid;
	wire branch_6_clk;
	wire branch_6_rst;
	wire [31 : 0] branch_6_in1_data;
	wire branch_6_in1_ready;
	wire branch_6_in1_valid;
	wire branch_6_in2_data;
	wire branch_6_in2_ready;
	wire branch_6_in2_valid;
	wire [31 : 0] branch_6_out1_data;
	wire branch_6_out1_ready;
	wire branch_6_out1_valid;
	wire [31 : 0] branch_6_out2_data;
	wire branch_6_out2_ready;
	wire branch_6_out2_valid;
	wire fork_30_clk;
	wire fork_30_rst;
	wire fork_30_in1_data;
	wire fork_30_in1_ready;
	wire fork_30_in1_valid;
	wire fork_30_out1_data;
	wire fork_30_out1_ready;
	wire fork_30_out1_valid;
	wire fork_30_out2_data;
	wire fork_30_out2_ready;
	wire fork_30_out2_valid;
	wire fork_30_out3_data;
	wire fork_30_out3_ready;
	wire fork_30_out3_valid;
	wire fork_30_out4_data;
	wire fork_30_out4_ready;
	wire fork_30_out4_valid;
	wire fork_30_out5_data;
	wire fork_30_out5_ready;
	wire fork_30_out5_valid;
	wire branch_7_clk;
	wire branch_7_rst;
	wire [5 : 0] branch_7_in1_data;
	wire branch_7_in1_ready;
	wire branch_7_in1_valid;
	wire branch_7_in2_data;
	wire branch_7_in2_ready;
	wire branch_7_in2_valid;
	wire [5 : 0] branch_7_out1_data;
	wire branch_7_out1_ready;
	wire branch_7_out1_valid;
	wire [5 : 0] branch_7_out2_data;
	wire branch_7_out2_ready;
	wire branch_7_out2_valid;
	wire branch_8_clk;
	wire branch_8_rst;
	wire [5 : 0] branch_8_in1_data;
	wire branch_8_in1_ready;
	wire branch_8_in1_valid;
	wire branch_8_in2_data;
	wire branch_8_in2_ready;
	wire branch_8_in2_valid;
	wire [5 : 0] branch_8_out1_data;
	wire branch_8_out1_ready;
	wire branch_8_out1_valid;
	wire [5 : 0] branch_8_out2_data;
	wire branch_8_out2_ready;
	wire branch_8_out2_valid;
	wire branch_9_clk;
	wire branch_9_rst;
	wire [31 : 0] branch_9_in1_data;
	wire branch_9_in1_ready;
	wire branch_9_in1_valid;
	wire branch_9_in2_data;
	wire branch_9_in2_ready;
	wire branch_9_in2_valid;
	wire [31 : 0] branch_9_out1_data;
	wire branch_9_out1_ready;
	wire branch_9_out1_valid;
	wire [31 : 0] branch_9_out2_data;
	wire branch_9_out2_ready;
	wire branch_9_out2_valid;
	wire branch_10_clk;
	wire branch_10_rst;
	wire [31 : 0] branch_10_in1_data;
	wire branch_10_in1_ready;
	wire branch_10_in1_valid;
	wire branch_10_in2_data;
	wire branch_10_in2_ready;
	wire branch_10_in2_valid;
	wire [31 : 0] branch_10_out1_data;
	wire branch_10_out1_ready;
	wire branch_10_out1_valid;
	wire [31 : 0] branch_10_out2_data;
	wire branch_10_out2_ready;
	wire branch_10_out2_valid;
	wire fork_31_clk;
	wire fork_31_rst;
	wire fork_31_in1_data;
	wire fork_31_in1_ready;
	wire fork_31_in1_valid;
	wire fork_31_out1_data;
	wire fork_31_out1_ready;
	wire fork_31_out1_valid;
	wire fork_31_out2_data;
	wire fork_31_out2_ready;
	wire fork_31_out2_valid;
	wire fork_31_out3_data;
	wire fork_31_out3_ready;
	wire fork_31_out3_valid;
	wire fork_31_out4_data;
	wire fork_31_out4_ready;
	wire fork_31_out4_valid;
	wire fork_31_out5_data;
	wire fork_31_out5_ready;
	wire fork_31_out5_valid;
	wire branch_11_clk;
	wire branch_11_rst;
	wire [5 : 0] branch_11_in1_data;
	wire branch_11_in1_ready;
	wire branch_11_in1_valid;
	wire branch_11_in2_data;
	wire branch_11_in2_ready;
	wire branch_11_in2_valid;
	wire [5 : 0] branch_11_out1_data;
	wire branch_11_out1_ready;
	wire branch_11_out1_valid;
	wire [5 : 0] branch_11_out2_data;
	wire branch_11_out2_ready;
	wire branch_11_out2_valid;
	wire branch_12_clk;
	wire branch_12_rst;
	wire [31 : 0] branch_12_in1_data;
	wire branch_12_in1_ready;
	wire branch_12_in1_valid;
	wire branch_12_in2_data;
	wire branch_12_in2_ready;
	wire branch_12_in2_valid;
	wire [31 : 0] branch_12_out1_data;
	wire branch_12_out1_ready;
	wire branch_12_out1_valid;
	wire [31 : 0] branch_12_out2_data;
	wire branch_12_out2_ready;
	wire branch_12_out2_valid;
	wire branch_13_clk;
	wire branch_13_rst;
	wire [31 : 0] branch_13_in1_data;
	wire branch_13_in1_ready;
	wire branch_13_in1_valid;
	wire branch_13_in2_data;
	wire branch_13_in2_ready;
	wire branch_13_in2_valid;
	wire [31 : 0] branch_13_out1_data;
	wire branch_13_out1_ready;
	wire branch_13_out1_valid;
	wire [31 : 0] branch_13_out2_data;
	wire branch_13_out2_ready;
	wire branch_13_out2_valid;
	wire fork_32_clk;
	wire fork_32_rst;
	wire fork_32_in1_data;
	wire fork_32_in1_ready;
	wire fork_32_in1_valid;
	wire fork_32_out1_data;
	wire fork_32_out1_ready;
	wire fork_32_out1_valid;
	wire fork_32_out2_data;
	wire fork_32_out2_ready;
	wire fork_32_out2_valid;
	wire fork_32_out3_data;
	wire fork_32_out3_ready;
	wire fork_32_out3_valid;
	wire fork_32_out4_data;
	wire fork_32_out4_ready;
	wire fork_32_out4_valid;
	wire branch_14_clk;
	wire branch_14_rst;
	wire branch_14_in1_data;
	wire branch_14_in1_ready;
	wire branch_14_in1_valid;
	wire branch_14_in2_data;
	wire branch_14_in2_ready;
	wire branch_14_in2_valid;
	wire branch_14_out1_data;
	wire branch_14_out1_ready;
	wire branch_14_out1_valid;
	wire branch_14_out2_data;
	wire branch_14_out2_ready;
	wire branch_14_out2_valid;
	wire branch_15_clk;
	wire branch_15_rst;
	wire [31 : 0] branch_15_in1_data;
	wire branch_15_in1_ready;
	wire branch_15_in1_valid;
	wire branch_15_in2_data;
	wire branch_15_in2_ready;
	wire branch_15_in2_valid;
	wire [31 : 0] branch_15_out1_data;
	wire branch_15_out1_ready;
	wire branch_15_out1_valid;
	wire [31 : 0] branch_15_out2_data;
	wire branch_15_out2_ready;
	wire branch_15_out2_valid;
	wire branch_16_clk;
	wire branch_16_rst;
	wire [31 : 0] branch_16_in1_data;
	wire branch_16_in1_ready;
	wire branch_16_in1_valid;
	wire branch_16_in2_data;
	wire branch_16_in2_ready;
	wire branch_16_in2_valid;
	wire [31 : 0] branch_16_out1_data;
	wire branch_16_out1_ready;
	wire branch_16_out1_valid;
	wire [31 : 0] branch_16_out2_data;
	wire branch_16_out2_ready;
	wire branch_16_out2_valid;
	wire fork_33_clk;
	wire fork_33_rst;
	wire fork_33_in1_data;
	wire fork_33_in1_ready;
	wire fork_33_in1_valid;
	wire fork_33_out1_data;
	wire fork_33_out1_ready;
	wire fork_33_out1_valid;
	wire fork_33_out2_data;
	wire fork_33_out2_ready;
	wire fork_33_out2_valid;
	wire fork_33_out3_data;
	wire fork_33_out3_ready;
	wire fork_33_out3_valid;
	wire fork_33_out4_data;
	wire fork_33_out4_ready;
	wire fork_33_out4_valid;
	wire branch_17_clk;
	wire branch_17_rst;
	wire [31 : 0] branch_17_in1_data;
	wire branch_17_in1_ready;
	wire branch_17_in1_valid;
	wire branch_17_in2_data;
	wire branch_17_in2_ready;
	wire branch_17_in2_valid;
	wire [31 : 0] branch_17_out1_data;
	wire branch_17_out1_ready;
	wire branch_17_out1_valid;
	wire [31 : 0] branch_17_out2_data;
	wire branch_17_out2_ready;
	wire branch_17_out2_valid;
	wire branch_18_clk;
	wire branch_18_rst;
	wire branch_18_in1_data;
	wire branch_18_in1_ready;
	wire branch_18_in1_valid;
	wire branch_18_in2_data;
	wire branch_18_in2_ready;
	wire branch_18_in2_valid;
	wire branch_18_out1_data;
	wire branch_18_out1_ready;
	wire branch_18_out1_valid;
	wire branch_18_out2_data;
	wire branch_18_out2_ready;
	wire branch_18_out2_valid;
	wire branch_19_clk;
	wire branch_19_rst;
	wire [31 : 0] branch_19_in1_data;
	wire branch_19_in1_ready;
	wire branch_19_in1_valid;
	wire branch_19_in2_data;
	wire branch_19_in2_ready;
	wire branch_19_in2_valid;
	wire [31 : 0] branch_19_out1_data;
	wire branch_19_out1_ready;
	wire branch_19_out1_valid;
	wire [31 : 0] branch_19_out2_data;
	wire branch_19_out2_ready;
	wire branch_19_out2_valid;
	wire branch_20_clk;
	wire branch_20_rst;
	wire [31 : 0] branch_20_in1_data;
	wire branch_20_in1_ready;
	wire branch_20_in1_valid;
	wire branch_20_in2_data;
	wire branch_20_in2_ready;
	wire branch_20_in2_valid;
	wire [31 : 0] branch_20_out1_data;
	wire branch_20_out1_ready;
	wire branch_20_out1_valid;
	wire [31 : 0] branch_20_out2_data;
	wire branch_20_out2_ready;
	wire branch_20_out2_valid;
	wire branch_21_clk;
	wire branch_21_rst;
	wire [5 : 0] branch_21_in1_data;
	wire branch_21_in1_ready;
	wire branch_21_in1_valid;
	wire branch_21_in2_data;
	wire branch_21_in2_ready;
	wire branch_21_in2_valid;
	wire [5 : 0] branch_21_out1_data;
	wire branch_21_out1_ready;
	wire branch_21_out1_valid;
	wire [5 : 0] branch_21_out2_data;
	wire branch_21_out2_ready;
	wire branch_21_out2_valid;
	wire fork_34_clk;
	wire fork_34_rst;
	wire fork_34_in1_data;
	wire fork_34_in1_ready;
	wire fork_34_in1_valid;
	wire fork_34_out1_data;
	wire fork_34_out1_ready;
	wire fork_34_out1_valid;
	wire fork_34_out2_data;
	wire fork_34_out2_ready;
	wire fork_34_out2_valid;
	wire fork_34_out3_data;
	wire fork_34_out3_ready;
	wire fork_34_out3_valid;
	wire fork_34_out4_data;
	wire fork_34_out4_ready;
	wire fork_34_out4_valid;
	wire fork_34_out5_data;
	wire fork_34_out5_ready;
	wire fork_34_out5_valid;
	wire fork_34_out6_data;
	wire fork_34_out6_ready;
	wire fork_34_out6_valid;
	wire branch_22_clk;
	wire branch_22_rst;
	wire [31 : 0] branch_22_in1_data;
	wire branch_22_in1_ready;
	wire branch_22_in1_valid;
	wire branch_22_in2_data;
	wire branch_22_in2_ready;
	wire branch_22_in2_valid;
	wire [31 : 0] branch_22_out1_data;
	wire branch_22_out1_ready;
	wire branch_22_out1_valid;
	wire [31 : 0] branch_22_out2_data;
	wire branch_22_out2_ready;
	wire branch_22_out2_valid;
	wire branch_23_clk;
	wire branch_23_rst;
	wire [5 : 0] branch_23_in1_data;
	wire branch_23_in1_ready;
	wire branch_23_in1_valid;
	wire branch_23_in2_data;
	wire branch_23_in2_ready;
	wire branch_23_in2_valid;
	wire [5 : 0] branch_23_out1_data;
	wire branch_23_out1_ready;
	wire branch_23_out1_valid;
	wire [5 : 0] branch_23_out2_data;
	wire branch_23_out2_ready;
	wire branch_23_out2_valid;
	wire branch_24_clk;
	wire branch_24_rst;
	wire [5 : 0] branch_24_in1_data;
	wire branch_24_in1_ready;
	wire branch_24_in1_valid;
	wire branch_24_in2_data;
	wire branch_24_in2_ready;
	wire branch_24_in2_valid;
	wire [5 : 0] branch_24_out1_data;
	wire branch_24_out1_ready;
	wire branch_24_out1_valid;
	wire [5 : 0] branch_24_out2_data;
	wire branch_24_out2_ready;
	wire branch_24_out2_valid;
	wire branch_25_clk;
	wire branch_25_rst;
	wire [31 : 0] branch_25_in1_data;
	wire branch_25_in1_ready;
	wire branch_25_in1_valid;
	wire branch_25_in2_data;
	wire branch_25_in2_ready;
	wire branch_25_in2_valid;
	wire [31 : 0] branch_25_out1_data;
	wire branch_25_out1_ready;
	wire branch_25_out1_valid;
	wire [31 : 0] branch_25_out2_data;
	wire branch_25_out2_ready;
	wire branch_25_out2_valid;
	wire branch_26_clk;
	wire branch_26_rst;
	wire [31 : 0] branch_26_in1_data;
	wire branch_26_in1_ready;
	wire branch_26_in1_valid;
	wire branch_26_in2_data;
	wire branch_26_in2_ready;
	wire branch_26_in2_valid;
	wire [31 : 0] branch_26_out1_data;
	wire branch_26_out1_ready;
	wire branch_26_out1_valid;
	wire [31 : 0] branch_26_out2_data;
	wire branch_26_out2_ready;
	wire branch_26_out2_valid;
	wire fork_35_clk;
	wire fork_35_rst;
	wire fork_35_in1_data;
	wire fork_35_in1_ready;
	wire fork_35_in1_valid;
	wire fork_35_out1_data;
	wire fork_35_out1_ready;
	wire fork_35_out1_valid;
	wire fork_35_out2_data;
	wire fork_35_out2_ready;
	wire fork_35_out2_valid;
	wire fork_35_out3_data;
	wire fork_35_out3_ready;
	wire fork_35_out3_valid;
	wire fork_35_out4_data;
	wire fork_35_out4_ready;
	wire fork_35_out4_valid;
	wire fork_35_out5_data;
	wire fork_35_out5_ready;
	wire fork_35_out5_valid;
	wire fork_35_out6_data;
	wire fork_35_out6_ready;
	wire fork_35_out6_valid;
	wire branch_27_clk;
	wire branch_27_rst;
	wire [31 : 0] branch_27_in1_data;
	wire branch_27_in1_ready;
	wire branch_27_in1_valid;
	wire branch_27_in2_data;
	wire branch_27_in2_ready;
	wire branch_27_in2_valid;
	wire [31 : 0] branch_27_out1_data;
	wire branch_27_out1_ready;
	wire branch_27_out1_valid;
	wire [31 : 0] branch_27_out2_data;
	wire branch_27_out2_ready;
	wire branch_27_out2_valid;
	wire branch_28_clk;
	wire branch_28_rst;
	wire [5 : 0] branch_28_in1_data;
	wire branch_28_in1_ready;
	wire branch_28_in1_valid;
	wire branch_28_in2_data;
	wire branch_28_in2_ready;
	wire branch_28_in2_valid;
	wire [5 : 0] branch_28_out1_data;
	wire branch_28_out1_ready;
	wire branch_28_out1_valid;
	wire [5 : 0] branch_28_out2_data;
	wire branch_28_out2_ready;
	wire branch_28_out2_valid;
	wire branch_29_clk;
	wire branch_29_rst;
	wire [31 : 0] branch_29_in1_data;
	wire branch_29_in1_ready;
	wire branch_29_in1_valid;
	wire branch_29_in2_data;
	wire branch_29_in2_ready;
	wire branch_29_in2_valid;
	wire [31 : 0] branch_29_out1_data;
	wire branch_29_out1_ready;
	wire branch_29_out1_valid;
	wire [31 : 0] branch_29_out2_data;
	wire branch_29_out2_ready;
	wire branch_29_out2_valid;
	wire fork_36_clk;
	wire fork_36_rst;
	wire fork_36_in1_data;
	wire fork_36_in1_ready;
	wire fork_36_in1_valid;
	wire fork_36_out1_data;
	wire fork_36_out1_ready;
	wire fork_36_out1_valid;
	wire fork_36_out2_data;
	wire fork_36_out2_ready;
	wire fork_36_out2_valid;
	wire fork_36_out3_data;
	wire fork_36_out3_ready;
	wire fork_36_out3_valid;
	wire fork_36_out4_data;
	wire fork_36_out4_ready;
	wire fork_36_out4_valid;
	wire branch_30_clk;
	wire branch_30_rst;
	wire branch_30_in1_data;
	wire branch_30_in1_ready;
	wire branch_30_in1_valid;
	wire branch_30_in2_data;
	wire branch_30_in2_ready;
	wire branch_30_in2_valid;
	wire branch_30_out1_data;
	wire branch_30_out1_ready;
	wire branch_30_out1_valid;
	wire branch_30_out2_data;
	wire branch_30_out2_ready;
	wire branch_30_out2_valid;
	wire branch_31_clk;
	wire branch_31_rst;
	wire [31 : 0] branch_31_in1_data;
	wire branch_31_in1_ready;
	wire branch_31_in1_valid;
	wire branch_31_in2_data;
	wire branch_31_in2_ready;
	wire branch_31_in2_valid;
	wire [31 : 0] branch_31_out1_data;
	wire branch_31_out1_ready;
	wire branch_31_out1_valid;
	wire [31 : 0] branch_31_out2_data;
	wire branch_31_out2_ready;
	wire branch_31_out2_valid;
	wire fork_37_clk;
	wire fork_37_rst;
	wire fork_37_in1_data;
	wire fork_37_in1_ready;
	wire fork_37_in1_valid;
	wire fork_37_out1_data;
	wire fork_37_out1_ready;
	wire fork_37_out1_valid;
	wire fork_37_out2_data;
	wire fork_37_out2_ready;
	wire fork_37_out2_valid;
	wire fork_37_out3_data;
	wire fork_37_out3_ready;
	wire fork_37_out3_valid;
	wire branch_32_clk;
	wire branch_32_rst;
	wire [5 : 0] branch_32_in1_data;
	wire branch_32_in1_ready;
	wire branch_32_in1_valid;
	wire branch_32_in2_data;
	wire branch_32_in2_ready;
	wire branch_32_in2_valid;
	wire [5 : 0] branch_32_out1_data;
	wire branch_32_out1_ready;
	wire branch_32_out1_valid;
	wire [5 : 0] branch_32_out2_data;
	wire branch_32_out2_ready;
	wire branch_32_out2_valid;
	wire branch_33_clk;
	wire branch_33_rst;
	wire [31 : 0] branch_33_in1_data;
	wire branch_33_in1_ready;
	wire branch_33_in1_valid;
	wire branch_33_in2_data;
	wire branch_33_in2_ready;
	wire branch_33_in2_valid;
	wire [31 : 0] branch_33_out1_data;
	wire branch_33_out1_ready;
	wire branch_33_out1_valid;
	wire [31 : 0] branch_33_out2_data;
	wire branch_33_out2_ready;
	wire branch_33_out2_valid;
	wire fork_38_clk;
	wire fork_38_rst;
	wire fork_38_in1_data;
	wire fork_38_in1_ready;
	wire fork_38_in1_valid;
	wire fork_38_out1_data;
	wire fork_38_out1_ready;
	wire fork_38_out1_valid;
	wire fork_38_out2_data;
	wire fork_38_out2_ready;
	wire fork_38_out2_valid;
	wire fork_38_out3_data;
	wire fork_38_out3_ready;
	wire fork_38_out3_valid;
	wire branch_34_clk;
	wire branch_34_rst;
	wire branch_34_in1_data;
	wire branch_34_in1_ready;
	wire branch_34_in1_valid;
	wire branch_34_in2_data;
	wire branch_34_in2_ready;
	wire branch_34_in2_valid;
	wire branch_34_out1_data;
	wire branch_34_out1_ready;
	wire branch_34_out1_valid;
	wire branch_34_out2_data;
	wire branch_34_out2_ready;
	wire branch_34_out2_valid;
	wire branch_35_clk;
	wire branch_35_rst;
	wire [31 : 0] branch_35_in1_data;
	wire branch_35_in1_ready;
	wire branch_35_in1_valid;
	wire branch_35_in2_data;
	wire branch_35_in2_ready;
	wire branch_35_in2_valid;
	wire [31 : 0] branch_35_out1_data;
	wire branch_35_out1_ready;
	wire branch_35_out1_valid;
	wire [31 : 0] branch_35_out2_data;
	wire branch_35_out2_ready;
	wire branch_35_out2_valid;
	wire fork_39_clk;
	wire fork_39_rst;
	wire fork_39_in1_data;
	wire fork_39_in1_ready;
	wire fork_39_in1_valid;
	wire fork_39_out1_data;
	wire fork_39_out1_ready;
	wire fork_39_out1_valid;
	wire fork_39_out2_data;
	wire fork_39_out2_ready;
	wire fork_39_out2_valid;
	wire fork_39_out3_data;
	wire fork_39_out3_ready;
	wire fork_39_out3_valid;
	wire branch_36_clk;
	wire branch_36_rst;
	wire [31 : 0] branch_36_in1_data;
	wire branch_36_in1_ready;
	wire branch_36_in1_valid;
	wire branch_36_in2_data;
	wire branch_36_in2_ready;
	wire branch_36_in2_valid;
	wire [31 : 0] branch_36_out1_data;
	wire branch_36_out1_ready;
	wire branch_36_out1_valid;
	wire [31 : 0] branch_36_out2_data;
	wire branch_36_out2_ready;
	wire branch_36_out2_valid;
	wire branch_37_clk;
	wire branch_37_rst;
	wire branch_37_in1_data;
	wire branch_37_in1_ready;
	wire branch_37_in1_valid;
	wire branch_37_in2_data;
	wire branch_37_in2_ready;
	wire branch_37_in2_valid;
	wire branch_37_out1_data;
	wire branch_37_out1_ready;
	wire branch_37_out1_valid;
	wire branch_37_out2_data;
	wire branch_37_out2_ready;
	wire branch_37_out2_valid;
	wire branch_38_clk;
	wire branch_38_rst;
	wire [31 : 0] branch_38_in1_data;
	wire branch_38_in1_ready;
	wire branch_38_in1_valid;
	wire branch_38_in2_data;
	wire branch_38_in2_ready;
	wire branch_38_in2_valid;
	wire [31 : 0] branch_38_out1_data;
	wire branch_38_out1_ready;
	wire branch_38_out1_valid;
	wire [31 : 0] branch_38_out2_data;
	wire branch_38_out2_ready;
	wire branch_38_out2_valid;
	wire branch_39_clk;
	wire branch_39_rst;
	wire [5 : 0] branch_39_in1_data;
	wire branch_39_in1_ready;
	wire branch_39_in1_valid;
	wire branch_39_in2_data;
	wire branch_39_in2_ready;
	wire branch_39_in2_valid;
	wire [5 : 0] branch_39_out1_data;
	wire branch_39_out1_ready;
	wire branch_39_out1_valid;
	wire [5 : 0] branch_39_out2_data;
	wire branch_39_out2_ready;
	wire branch_39_out2_valid;
	wire fork_40_clk;
	wire fork_40_rst;
	wire fork_40_in1_data;
	wire fork_40_in1_ready;
	wire fork_40_in1_valid;
	wire fork_40_out1_data;
	wire fork_40_out1_ready;
	wire fork_40_out1_valid;
	wire fork_40_out2_data;
	wire fork_40_out2_ready;
	wire fork_40_out2_valid;
	wire fork_40_out3_data;
	wire fork_40_out3_ready;
	wire fork_40_out3_valid;
	wire fork_40_out4_data;
	wire fork_40_out4_ready;
	wire fork_40_out4_valid;
	wire fork_40_out5_data;
	wire fork_40_out5_ready;
	wire fork_40_out5_valid;
	wire branch_40_clk;
	wire branch_40_rst;
	wire [31 : 0] branch_40_in1_data;
	wire branch_40_in1_ready;
	wire branch_40_in1_valid;
	wire branch_40_in2_data;
	wire branch_40_in2_ready;
	wire branch_40_in2_valid;
	wire [31 : 0] branch_40_out1_data;
	wire branch_40_out1_ready;
	wire branch_40_out1_valid;
	wire [31 : 0] branch_40_out2_data;
	wire branch_40_out2_ready;
	wire branch_40_out2_valid;
	wire branch_41_clk;
	wire branch_41_rst;
	wire [5 : 0] branch_41_in1_data;
	wire branch_41_in1_ready;
	wire branch_41_in1_valid;
	wire branch_41_in2_data;
	wire branch_41_in2_ready;
	wire branch_41_in2_valid;
	wire [5 : 0] branch_41_out1_data;
	wire branch_41_out1_ready;
	wire branch_41_out1_valid;
	wire [5 : 0] branch_41_out2_data;
	wire branch_41_out2_ready;
	wire branch_41_out2_valid;
	wire branch_42_clk;
	wire branch_42_rst;
	wire [5 : 0] branch_42_in1_data;
	wire branch_42_in1_ready;
	wire branch_42_in1_valid;
	wire branch_42_in2_data;
	wire branch_42_in2_ready;
	wire branch_42_in2_valid;
	wire [5 : 0] branch_42_out1_data;
	wire branch_42_out1_ready;
	wire branch_42_out1_valid;
	wire [5 : 0] branch_42_out2_data;
	wire branch_42_out2_ready;
	wire branch_42_out2_valid;
	wire branch_43_clk;
	wire branch_43_rst;
	wire [31 : 0] branch_43_in1_data;
	wire branch_43_in1_ready;
	wire branch_43_in1_valid;
	wire branch_43_in2_data;
	wire branch_43_in2_ready;
	wire branch_43_in2_valid;
	wire [31 : 0] branch_43_out1_data;
	wire branch_43_out1_ready;
	wire branch_43_out1_valid;
	wire [31 : 0] branch_43_out2_data;
	wire branch_43_out2_ready;
	wire branch_43_out2_valid;
	wire fork_41_clk;
	wire fork_41_rst;
	wire fork_41_in1_data;
	wire fork_41_in1_ready;
	wire fork_41_in1_valid;
	wire fork_41_out1_data;
	wire fork_41_out1_ready;
	wire fork_41_out1_valid;
	wire fork_41_out2_data;
	wire fork_41_out2_ready;
	wire fork_41_out2_valid;
	wire fork_41_out3_data;
	wire fork_41_out3_ready;
	wire fork_41_out3_valid;
	wire fork_41_out4_data;
	wire fork_41_out4_ready;
	wire fork_41_out4_valid;
	wire fork_41_out5_data;
	wire fork_41_out5_ready;
	wire fork_41_out5_valid;
	wire branch_44_clk;
	wire branch_44_rst;
	wire [31 : 0] branch_44_in1_data;
	wire branch_44_in1_ready;
	wire branch_44_in1_valid;
	wire branch_44_in2_data;
	wire branch_44_in2_ready;
	wire branch_44_in2_valid;
	wire [31 : 0] branch_44_out1_data;
	wire branch_44_out1_ready;
	wire branch_44_out1_valid;
	wire [31 : 0] branch_44_out2_data;
	wire branch_44_out2_ready;
	wire branch_44_out2_valid;
	wire branch_45_clk;
	wire branch_45_rst;
	wire [5 : 0] branch_45_in1_data;
	wire branch_45_in1_ready;
	wire branch_45_in1_valid;
	wire branch_45_in2_data;
	wire branch_45_in2_ready;
	wire branch_45_in2_valid;
	wire [5 : 0] branch_45_out1_data;
	wire branch_45_out1_ready;
	wire branch_45_out1_valid;
	wire [5 : 0] branch_45_out2_data;
	wire branch_45_out2_ready;
	wire branch_45_out2_valid;
	wire fork_42_clk;
	wire fork_42_rst;
	wire fork_42_in1_data;
	wire fork_42_in1_ready;
	wire fork_42_in1_valid;
	wire fork_42_out1_data;
	wire fork_42_out1_ready;
	wire fork_42_out1_valid;
	wire fork_42_out2_data;
	wire fork_42_out2_ready;
	wire fork_42_out2_valid;
	wire fork_42_out3_data;
	wire fork_42_out3_ready;
	wire fork_42_out3_valid;
	wire MC_A_clk;
	wire MC_A_rst;
	wire [31 : 0] MC_A_in1_data;
	wire MC_A_in1_ready;
	wire MC_A_in1_valid;
	wire [11 : 0] MC_A_in2_data;
	wire MC_A_in2_ready;
	wire MC_A_in2_valid;
	wire [11 : 0] MC_A_in3_data;
	wire MC_A_in3_ready;
	wire MC_A_in3_valid;
	wire [31 : 0] MC_A_in4_data;
	wire MC_A_in4_ready;
	wire MC_A_in4_valid;
	wire [11 : 0] MC_A_in5_data;
	wire MC_A_in5_ready;
	wire MC_A_in5_valid;
	wire [11 : 0] MC_A_in6_data;
	wire MC_A_in6_ready;
	wire MC_A_in6_valid;
	wire [31 : 0] MC_A_out1_data;
	wire MC_A_out1_ready;
	wire MC_A_out1_valid;
	wire [31 : 0] MC_A_out2_data;
	wire MC_A_out2_ready;
	wire MC_A_out2_valid;
	wire [31 : 0] MC_A_out3_data;
	wire MC_A_out3_ready;
	wire MC_A_out3_valid;
	wire MC_A_out4_data;
	wire MC_A_out4_ready;
	wire MC_A_out4_valid;
	wire MC_u1_clk;
	wire MC_u1_rst;
	wire [5 : 0] MC_u1_in1_data;
	wire MC_u1_in1_ready;
	wire MC_u1_in1_valid;
	wire [31 : 0] MC_u1_in2_data;
	wire MC_u1_in2_ready;
	wire MC_u1_in2_valid;
	wire [5 : 0] MC_u1_in3_data;
	wire MC_u1_in3_ready;
	wire MC_u1_in3_valid;
	wire [31 : 0] MC_u1_in4_data;
	wire MC_u1_in4_ready;
	wire MC_u1_in4_valid;
	wire [31 : 0] MC_u1_out1_data;
	wire MC_u1_out1_ready;
	wire MC_u1_out1_valid;
	wire MC_u1_out2_data;
	wire MC_u1_out2_ready;
	wire MC_u1_out2_valid;
	wire MC_v1_clk;
	wire MC_v1_rst;
	wire [5 : 0] MC_v1_in1_data;
	wire MC_v1_in1_ready;
	wire MC_v1_in1_valid;
	wire [31 : 0] MC_v1_in2_data;
	wire MC_v1_in2_ready;
	wire MC_v1_in2_valid;
	wire [5 : 0] MC_v1_in3_data;
	wire MC_v1_in3_ready;
	wire MC_v1_in3_valid;
	wire [31 : 0] MC_v1_in4_data;
	wire MC_v1_in4_ready;
	wire MC_v1_in4_valid;
	wire [31 : 0] MC_v1_out1_data;
	wire MC_v1_out1_ready;
	wire MC_v1_out1_valid;
	wire MC_v1_out2_data;
	wire MC_v1_out2_ready;
	wire MC_v1_out2_valid;
	wire MC_u2_clk;
	wire MC_u2_rst;
	wire [5 : 0] MC_u2_in1_data;
	wire MC_u2_in1_ready;
	wire MC_u2_in1_valid;
	wire [31 : 0] MC_u2_in2_data;
	wire MC_u2_in2_ready;
	wire MC_u2_in2_valid;
	wire [5 : 0] MC_u2_in3_data;
	wire MC_u2_in3_ready;
	wire MC_u2_in3_valid;
	wire [31 : 0] MC_u2_in4_data;
	wire MC_u2_in4_ready;
	wire MC_u2_in4_valid;
	wire [31 : 0] MC_u2_out1_data;
	wire MC_u2_out1_ready;
	wire MC_u2_out1_valid;
	wire MC_u2_out2_data;
	wire MC_u2_out2_ready;
	wire MC_u2_out2_valid;
	wire MC_v2_clk;
	wire MC_v2_rst;
	wire [5 : 0] MC_v2_in1_data;
	wire MC_v2_in1_ready;
	wire MC_v2_in1_valid;
	wire [31 : 0] MC_v2_in2_data;
	wire MC_v2_in2_ready;
	wire MC_v2_in2_valid;
	wire [5 : 0] MC_v2_in3_data;
	wire MC_v2_in3_ready;
	wire MC_v2_in3_valid;
	wire [31 : 0] MC_v2_in4_data;
	wire MC_v2_in4_ready;
	wire MC_v2_in4_valid;
	wire [31 : 0] MC_v2_out1_data;
	wire MC_v2_out1_ready;
	wire MC_v2_out1_valid;
	wire MC_v2_out2_data;
	wire MC_v2_out2_ready;
	wire MC_v2_out2_valid;
	wire cst_25_clk;
	wire cst_25_rst;
	wire cst_25_in1_data;
	wire cst_25_in1_ready;
	wire cst_25_in1_valid;
	wire cst_25_out1_data;
	wire cst_25_out1_ready;
	wire cst_25_out1_valid;
	wire MC_x_clk;
	wire MC_x_rst;
	wire [31 : 0] MC_x_in1_data;
	wire MC_x_in1_ready;
	wire MC_x_in1_valid;
	wire [31 : 0] MC_x_in2_data;
	wire MC_x_in2_ready;
	wire MC_x_in2_valid;
	wire [5 : 0] MC_x_in3_data;
	wire MC_x_in3_ready;
	wire MC_x_in3_valid;
	wire [5 : 0] MC_x_in4_data;
	wire MC_x_in4_ready;
	wire MC_x_in4_valid;
	wire [31 : 0] MC_x_in5_data;
	wire MC_x_in5_ready;
	wire MC_x_in5_valid;
	wire [5 : 0] MC_x_in6_data;
	wire MC_x_in6_ready;
	wire MC_x_in6_valid;
	wire [5 : 0] MC_x_in7_data;
	wire MC_x_in7_ready;
	wire MC_x_in7_valid;
	wire [31 : 0] MC_x_in8_data;
	wire MC_x_in8_ready;
	wire MC_x_in8_valid;
	wire [5 : 0] MC_x_in9_data;
	wire MC_x_in9_ready;
	wire MC_x_in9_valid;
	wire [31 : 0] MC_x_out1_data;
	wire MC_x_out1_ready;
	wire MC_x_out1_valid;
	wire [31 : 0] MC_x_out2_data;
	wire MC_x_out2_ready;
	wire MC_x_out2_valid;
	wire [31 : 0] MC_x_out3_data;
	wire MC_x_out3_ready;
	wire MC_x_out3_valid;
	wire MC_x_out4_data;
	wire MC_x_out4_ready;
	wire MC_x_out4_valid;
	wire MC_y_clk;
	wire MC_y_rst;
	wire [5 : 0] MC_y_in1_data;
	wire MC_y_in1_ready;
	wire MC_y_in1_valid;
	wire [31 : 0] MC_y_in2_data;
	wire MC_y_in2_ready;
	wire MC_y_in2_valid;
	wire [5 : 0] MC_y_in3_data;
	wire MC_y_in3_ready;
	wire MC_y_in3_valid;
	wire [31 : 0] MC_y_in4_data;
	wire MC_y_in4_ready;
	wire MC_y_in4_valid;
	wire [31 : 0] MC_y_out1_data;
	wire MC_y_out1_ready;
	wire MC_y_out1_valid;
	wire MC_y_out2_data;
	wire MC_y_out2_ready;
	wire MC_y_out2_valid;
	wire cst_26_clk;
	wire cst_26_rst;
	wire cst_26_in1_data;
	wire cst_26_in1_ready;
	wire cst_26_in1_valid;
	wire cst_26_out1_data;
	wire cst_26_out1_ready;
	wire cst_26_out1_valid;
	wire MC_z_clk;
	wire MC_z_rst;
	wire [5 : 0] MC_z_in1_data;
	wire MC_z_in1_ready;
	wire MC_z_in1_valid;
	wire [31 : 0] MC_z_in2_data;
	wire MC_z_in2_ready;
	wire MC_z_in2_valid;
	wire [5 : 0] MC_z_in3_data;
	wire MC_z_in3_ready;
	wire MC_z_in3_valid;
	wire [31 : 0] MC_z_in4_data;
	wire MC_z_in4_ready;
	wire MC_z_in4_valid;
	wire [31 : 0] MC_z_out1_data;
	wire MC_z_out1_ready;
	wire MC_z_out1_valid;
	wire MC_z_out2_data;
	wire MC_z_out2_ready;
	wire MC_z_out2_valid;
	wire cst_27_clk;
	wire cst_27_rst;
	wire cst_27_in1_data;
	wire cst_27_in1_ready;
	wire cst_27_in1_valid;
	wire cst_27_out1_data;
	wire cst_27_out1_ready;
	wire cst_27_out1_valid;
	wire MC_w_clk;
	wire MC_w_rst;
	wire [31 : 0] MC_w_in1_data;
	wire MC_w_in1_ready;
	wire MC_w_in1_valid;
	wire [5 : 0] MC_w_in2_data;
	wire MC_w_in2_ready;
	wire MC_w_in2_valid;
	wire [5 : 0] MC_w_in3_data;
	wire MC_w_in3_ready;
	wire MC_w_in3_valid;
	wire [31 : 0] MC_w_in4_data;
	wire MC_w_in4_ready;
	wire MC_w_in4_valid;
	wire [31 : 0] MC_w_out1_data;
	wire MC_w_out1_ready;
	wire MC_w_out1_valid;
	wire MC_w_out2_data;
	wire MC_w_out2_ready;
	wire MC_w_out2_valid;
	wire cst_28_clk;
	wire cst_28_rst;
	wire cst_28_in1_data;
	wire cst_28_in1_ready;
	wire cst_28_in1_valid;
	wire cst_28_out1_data;
	wire cst_28_out1_ready;
	wire cst_28_out1_valid;
	wire end_0_clk;
	wire end_0_rst;
	wire end_0_in1_data;
	wire end_0_in1_ready;
	wire end_0_in1_valid;
	wire end_0_in2_data;
	wire end_0_in2_ready;
	wire end_0_in2_valid;
	wire end_0_in3_data;
	wire end_0_in3_ready;
	wire end_0_in3_valid;
	wire end_0_in4_data;
	wire end_0_in4_ready;
	wire end_0_in4_valid;
	wire end_0_in5_data;
	wire end_0_in5_ready;
	wire end_0_in5_valid;
	wire end_0_in6_data;
	wire end_0_in6_ready;
	wire end_0_in6_valid;
	wire end_0_in7_data;
	wire end_0_in7_ready;
	wire end_0_in7_valid;
	wire end_0_in8_data;
	wire end_0_in8_ready;
	wire end_0_in8_valid;
	wire end_0_in9_data;
	wire end_0_in9_ready;
	wire end_0_in9_valid;
	wire end_0_in10_data;
	wire end_0_in10_ready;
	wire end_0_in10_valid;
	wire end_0_out1_data;
	wire end_0_out1_ready;
	wire end_0_out1_valid;
	wire start_0_clk;
	wire start_0_rst;
	wire start_0_in1_data;
	wire start_0_in1_ready;
	wire start_0_in1_valid;
	wire start_0_out1_data;
	wire start_0_out1_ready;
	wire start_0_out1_valid;
	wire forkC_44_clk;
	wire forkC_44_rst;
	wire forkC_44_in1_data;
	wire forkC_44_in1_ready;
	wire forkC_44_in1_valid;
	wire forkC_44_out1_data;
	wire forkC_44_out1_ready;
	wire forkC_44_out1_valid;
	wire forkC_44_out2_data;
	wire forkC_44_out2_ready;
	wire forkC_44_out2_valid;
	wire forkC_44_out3_data;
	wire forkC_44_out3_ready;
	wire forkC_44_out3_valid;
	wire branchC_46_clk;
	wire branchC_46_rst;
	wire branchC_46_in1_data;
	wire branchC_46_in1_ready;
	wire branchC_46_in1_valid;
	wire branchC_46_in2_data;
	wire branchC_46_in2_ready;
	wire branchC_46_in2_valid;
	wire branchC_46_out1_data;
	wire branchC_46_out1_ready;
	wire branchC_46_out1_valid;
	wire branchC_46_out2_data;
	wire branchC_46_out2_ready;
	wire branchC_46_out2_valid;
	wire phiC_28_clk;
	wire phiC_28_rst;
	wire phiC_28_in1_data;
	wire phiC_28_in1_ready;
	wire phiC_28_in1_valid;
	wire phiC_28_in2_data;
	wire phiC_28_in2_ready;
	wire phiC_28_in2_valid;
	wire phiC_28_out1_data;
	wire phiC_28_out1_ready;
	wire phiC_28_out1_valid;
	wire phiC_28_out2_data;
	wire phiC_28_out2_ready;
	wire phiC_28_out2_valid;
	wire forkC_45_clk;
	wire forkC_45_rst;
	wire forkC_45_in1_data;
	wire forkC_45_in1_ready;
	wire forkC_45_in1_valid;
	wire forkC_45_out1_data;
	wire forkC_45_out1_ready;
	wire forkC_45_out1_valid;
	wire forkC_45_out2_data;
	wire forkC_45_out2_ready;
	wire forkC_45_out2_valid;
	wire forkC_45_out3_data;
	wire forkC_45_out3_ready;
	wire forkC_45_out3_valid;
	wire branchC_47_clk;
	wire branchC_47_rst;
	wire branchC_47_in1_data;
	wire branchC_47_in1_ready;
	wire branchC_47_in1_valid;
	wire branchC_47_in2_data;
	wire branchC_47_in2_ready;
	wire branchC_47_in2_valid;
	wire branchC_47_out1_data;
	wire branchC_47_out1_ready;
	wire branchC_47_out1_valid;
	wire branchC_47_out2_data;
	wire branchC_47_out2_ready;
	wire branchC_47_out2_valid;
	wire phiC_29_clk;
	wire phiC_29_rst;
	wire phiC_29_in1_data;
	wire phiC_29_in1_ready;
	wire phiC_29_in1_valid;
	wire phiC_29_in2_data;
	wire phiC_29_in2_ready;
	wire phiC_29_in2_valid;
	wire phiC_29_out1_data;
	wire phiC_29_out1_ready;
	wire phiC_29_out1_valid;
	wire phiC_29_out2_data;
	wire phiC_29_out2_ready;
	wire phiC_29_out2_valid;
	wire forkC_46_clk;
	wire forkC_46_rst;
	wire forkC_46_in1_data;
	wire forkC_46_in1_ready;
	wire forkC_46_in1_valid;
	wire forkC_46_out1_data;
	wire forkC_46_out1_ready;
	wire forkC_46_out1_valid;
	wire forkC_46_out2_data;
	wire forkC_46_out2_ready;
	wire forkC_46_out2_valid;
	wire branchC_48_clk;
	wire branchC_48_rst;
	wire branchC_48_in1_data;
	wire branchC_48_in1_ready;
	wire branchC_48_in1_valid;
	wire branchC_48_in2_data;
	wire branchC_48_in2_ready;
	wire branchC_48_in2_valid;
	wire branchC_48_out1_data;
	wire branchC_48_out1_ready;
	wire branchC_48_out1_valid;
	wire branchC_48_out2_data;
	wire branchC_48_out2_ready;
	wire branchC_48_out2_valid;
	wire phiC_30_clk;
	wire phiC_30_rst;
	wire phiC_30_in1_data;
	wire phiC_30_in1_ready;
	wire phiC_30_in1_valid;
	wire phiC_30_out1_data;
	wire phiC_30_out1_ready;
	wire phiC_30_out1_valid;
	wire branchC_49_clk;
	wire branchC_49_rst;
	wire branchC_49_in1_data;
	wire branchC_49_in1_ready;
	wire branchC_49_in1_valid;
	wire branchC_49_in2_data;
	wire branchC_49_in2_ready;
	wire branchC_49_in2_valid;
	wire branchC_49_out1_data;
	wire branchC_49_out1_ready;
	wire branchC_49_out1_valid;
	wire branchC_49_out2_data;
	wire branchC_49_out2_ready;
	wire branchC_49_out2_valid;
	wire phiC_31_clk;
	wire phiC_31_rst;
	wire phiC_31_in1_data;
	wire phiC_31_in1_ready;
	wire phiC_31_in1_valid;
	wire phiC_31_out1_data;
	wire phiC_31_out1_ready;
	wire phiC_31_out1_valid;
	wire forkC_48_clk;
	wire forkC_48_rst;
	wire forkC_48_in1_data;
	wire forkC_48_in1_ready;
	wire forkC_48_in1_valid;
	wire forkC_48_out1_data;
	wire forkC_48_out1_ready;
	wire forkC_48_out1_valid;
	wire forkC_48_out2_data;
	wire forkC_48_out2_ready;
	wire forkC_48_out2_valid;
	wire forkC_48_out3_data;
	wire forkC_48_out3_ready;
	wire forkC_48_out3_valid;
	wire branchC_50_clk;
	wire branchC_50_rst;
	wire branchC_50_in1_data;
	wire branchC_50_in1_ready;
	wire branchC_50_in1_valid;
	wire branchC_50_in2_data;
	wire branchC_50_in2_ready;
	wire branchC_50_in2_valid;
	wire branchC_50_out1_data;
	wire branchC_50_out1_ready;
	wire branchC_50_out1_valid;
	wire branchC_50_out2_data;
	wire branchC_50_out2_ready;
	wire branchC_50_out2_valid;
	wire phiC_32_clk;
	wire phiC_32_rst;
	wire phiC_32_in1_data;
	wire phiC_32_in1_ready;
	wire phiC_32_in1_valid;
	wire phiC_32_in2_data;
	wire phiC_32_in2_ready;
	wire phiC_32_in2_valid;
	wire phiC_32_out1_data;
	wire phiC_32_out1_ready;
	wire phiC_32_out1_valid;
	wire phiC_32_out2_data;
	wire phiC_32_out2_ready;
	wire phiC_32_out2_valid;
	wire forkC_49_clk;
	wire forkC_49_rst;
	wire forkC_49_in1_data;
	wire forkC_49_in1_ready;
	wire forkC_49_in1_valid;
	wire forkC_49_out1_data;
	wire forkC_49_out1_ready;
	wire forkC_49_out1_valid;
	wire forkC_49_out2_data;
	wire forkC_49_out2_ready;
	wire forkC_49_out2_valid;
	wire forkC_49_out3_data;
	wire forkC_49_out3_ready;
	wire forkC_49_out3_valid;
	wire branchC_51_clk;
	wire branchC_51_rst;
	wire branchC_51_in1_data;
	wire branchC_51_in1_ready;
	wire branchC_51_in1_valid;
	wire branchC_51_in2_data;
	wire branchC_51_in2_ready;
	wire branchC_51_in2_valid;
	wire branchC_51_out1_data;
	wire branchC_51_out1_ready;
	wire branchC_51_out1_valid;
	wire branchC_51_out2_data;
	wire branchC_51_out2_ready;
	wire branchC_51_out2_valid;
	wire phiC_33_clk;
	wire phiC_33_rst;
	wire phiC_33_in1_data;
	wire phiC_33_in1_ready;
	wire phiC_33_in1_valid;
	wire phiC_33_in2_data;
	wire phiC_33_in2_ready;
	wire phiC_33_in2_valid;
	wire phiC_33_out1_data;
	wire phiC_33_out1_ready;
	wire phiC_33_out1_valid;
	wire phiC_33_out2_data;
	wire phiC_33_out2_ready;
	wire phiC_33_out2_valid;
	wire branchC_52_clk;
	wire branchC_52_rst;
	wire branchC_52_in1_data;
	wire branchC_52_in1_ready;
	wire branchC_52_in1_valid;
	wire branchC_52_in2_data;
	wire branchC_52_in2_ready;
	wire branchC_52_in2_valid;
	wire branchC_52_out1_data;
	wire branchC_52_out1_ready;
	wire branchC_52_out1_valid;
	wire branchC_52_out2_data;
	wire branchC_52_out2_ready;
	wire branchC_52_out2_valid;
	wire phiC_34_clk;
	wire phiC_34_rst;
	wire phiC_34_in1_data;
	wire phiC_34_in1_ready;
	wire phiC_34_in1_valid;
	wire phiC_34_out1_data;
	wire phiC_34_out1_ready;
	wire phiC_34_out1_valid;
	wire forkC_51_clk;
	wire forkC_51_rst;
	wire forkC_51_in1_data;
	wire forkC_51_in1_ready;
	wire forkC_51_in1_valid;
	wire forkC_51_out1_data;
	wire forkC_51_out1_ready;
	wire forkC_51_out1_valid;
	wire forkC_51_out2_data;
	wire forkC_51_out2_ready;
	wire forkC_51_out2_valid;
	wire branchC_53_clk;
	wire branchC_53_rst;
	wire branchC_53_in1_data;
	wire branchC_53_in1_ready;
	wire branchC_53_in1_valid;
	wire branchC_53_in2_data;
	wire branchC_53_in2_ready;
	wire branchC_53_in2_valid;
	wire branchC_53_out1_data;
	wire branchC_53_out1_ready;
	wire branchC_53_out1_valid;
	wire branchC_53_out2_data;
	wire branchC_53_out2_ready;
	wire branchC_53_out2_valid;
	wire phiC_35_clk;
	wire phiC_35_rst;
	wire phiC_35_in1_data;
	wire phiC_35_in1_ready;
	wire phiC_35_in1_valid;
	wire phiC_35_out1_data;
	wire phiC_35_out1_ready;
	wire phiC_35_out1_valid;
	wire forkC_52_clk;
	wire forkC_52_rst;
	wire forkC_52_in1_data;
	wire forkC_52_in1_ready;
	wire forkC_52_in1_valid;
	wire forkC_52_out1_data;
	wire forkC_52_out1_ready;
	wire forkC_52_out1_valid;
	wire forkC_52_out2_data;
	wire forkC_52_out2_ready;
	wire forkC_52_out2_valid;
	wire forkC_52_out3_data;
	wire forkC_52_out3_ready;
	wire forkC_52_out3_valid;
	wire branchC_54_clk;
	wire branchC_54_rst;
	wire branchC_54_in1_data;
	wire branchC_54_in1_ready;
	wire branchC_54_in1_valid;
	wire branchC_54_in2_data;
	wire branchC_54_in2_ready;
	wire branchC_54_in2_valid;
	wire branchC_54_out1_data;
	wire branchC_54_out1_ready;
	wire branchC_54_out1_valid;
	wire branchC_54_out2_data;
	wire branchC_54_out2_ready;
	wire branchC_54_out2_valid;
	wire phiC_36_clk;
	wire phiC_36_rst;
	wire phiC_36_in1_data;
	wire phiC_36_in1_ready;
	wire phiC_36_in1_valid;
	wire phiC_36_in2_data;
	wire phiC_36_in2_ready;
	wire phiC_36_in2_valid;
	wire phiC_36_out1_data;
	wire phiC_36_out1_ready;
	wire phiC_36_out1_valid;
	wire phiC_36_out2_data;
	wire phiC_36_out2_ready;
	wire phiC_36_out2_valid;
	wire forkC_53_clk;
	wire forkC_53_rst;
	wire forkC_53_in1_data;
	wire forkC_53_in1_ready;
	wire forkC_53_in1_valid;
	wire forkC_53_out1_data;
	wire forkC_53_out1_ready;
	wire forkC_53_out1_valid;
	wire forkC_53_out2_data;
	wire forkC_53_out2_ready;
	wire forkC_53_out2_valid;
	wire branchC_55_clk;
	wire branchC_55_rst;
	wire branchC_55_in1_data;
	wire branchC_55_in1_ready;
	wire branchC_55_in1_valid;
	wire branchC_55_in2_data;
	wire branchC_55_in2_ready;
	wire branchC_55_in2_valid;
	wire branchC_55_out1_data;
	wire branchC_55_out1_ready;
	wire branchC_55_out1_valid;
	wire branchC_55_out2_data;
	wire branchC_55_out2_ready;
	wire branchC_55_out2_valid;
	wire phiC_37_clk;
	wire phiC_37_rst;
	wire phiC_37_in1_data;
	wire phiC_37_in1_ready;
	wire phiC_37_in1_valid;
	wire phiC_37_out1_data;
	wire phiC_37_out1_ready;
	wire phiC_37_out1_valid;
	wire forkC_54_clk;
	wire forkC_54_rst;
	wire forkC_54_in1_data;
	wire forkC_54_in1_ready;
	wire forkC_54_in1_valid;
	wire forkC_54_out1_data;
	wire forkC_54_out1_ready;
	wire forkC_54_out1_valid;
	wire forkC_54_out2_data;
	wire forkC_54_out2_ready;
	wire forkC_54_out2_valid;
	wire forkC_54_out3_data;
	wire forkC_54_out3_ready;
	wire forkC_54_out3_valid;
	wire branchC_56_clk;
	wire branchC_56_rst;
	wire branchC_56_in1_data;
	wire branchC_56_in1_ready;
	wire branchC_56_in1_valid;
	wire branchC_56_in2_data;
	wire branchC_56_in2_ready;
	wire branchC_56_in2_valid;
	wire branchC_56_out1_data;
	wire branchC_56_out1_ready;
	wire branchC_56_out1_valid;
	wire branchC_56_out2_data;
	wire branchC_56_out2_ready;
	wire branchC_56_out2_valid;
	wire phiC_38_clk;
	wire phiC_38_rst;
	wire phiC_38_in1_data;
	wire phiC_38_in1_ready;
	wire phiC_38_in1_valid;
	wire phiC_38_in2_data;
	wire phiC_38_in2_ready;
	wire phiC_38_in2_valid;
	wire phiC_38_out1_data;
	wire phiC_38_out1_ready;
	wire phiC_38_out1_valid;
	wire phiC_38_out2_data;
	wire phiC_38_out2_ready;
	wire phiC_38_out2_valid;
	wire forkC_55_clk;
	wire forkC_55_rst;
	wire forkC_55_in1_data;
	wire forkC_55_in1_ready;
	wire forkC_55_in1_valid;
	wire forkC_55_out1_data;
	wire forkC_55_out1_ready;
	wire forkC_55_out1_valid;
	wire forkC_55_out2_data;
	wire forkC_55_out2_ready;
	wire forkC_55_out2_valid;
	wire forkC_55_out3_data;
	wire forkC_55_out3_ready;
	wire forkC_55_out3_valid;
	wire branchC_57_clk;
	wire branchC_57_rst;
	wire branchC_57_in1_data;
	wire branchC_57_in1_ready;
	wire branchC_57_in1_valid;
	wire branchC_57_in2_data;
	wire branchC_57_in2_ready;
	wire branchC_57_in2_valid;
	wire branchC_57_out1_data;
	wire branchC_57_out1_ready;
	wire branchC_57_out1_valid;
	wire branchC_57_out2_data;
	wire branchC_57_out2_ready;
	wire branchC_57_out2_valid;
	wire phiC_39_clk;
	wire phiC_39_rst;
	wire phiC_39_in1_data;
	wire phiC_39_in1_ready;
	wire phiC_39_in1_valid;
	wire phiC_39_in2_data;
	wire phiC_39_in2_ready;
	wire phiC_39_in2_valid;
	wire phiC_39_out1_data;
	wire phiC_39_out1_ready;
	wire phiC_39_out1_valid;
	wire phiC_39_out2_data;
	wire phiC_39_out2_ready;
	wire phiC_39_out2_valid;
	wire branchC_58_clk;
	wire branchC_58_rst;
	wire branchC_58_in1_data;
	wire branchC_58_in1_ready;
	wire branchC_58_in1_valid;
	wire branchC_58_in2_data;
	wire branchC_58_in2_ready;
	wire branchC_58_in2_valid;
	wire branchC_58_out1_data;
	wire branchC_58_out1_ready;
	wire branchC_58_out1_valid;
	wire branchC_58_out2_data;
	wire branchC_58_out2_ready;
	wire branchC_58_out2_valid;
	wire phiC_40_clk;
	wire phiC_40_rst;
	wire phiC_40_in1_data;
	wire phiC_40_in1_ready;
	wire phiC_40_in1_valid;
	wire phiC_40_out1_data;
	wire phiC_40_out1_ready;
	wire phiC_40_out1_valid;
	wire forkC_57_clk;
	wire forkC_57_rst;
	wire forkC_57_in1_data;
	wire forkC_57_in1_ready;
	wire forkC_57_in1_valid;
	wire forkC_57_out1_data;
	wire forkC_57_out1_ready;
	wire forkC_57_out1_valid;
	wire forkC_57_out2_data;
	wire forkC_57_out2_ready;
	wire forkC_57_out2_valid;
	wire branchC_59_clk;
	wire branchC_59_rst;
	wire branchC_59_in1_data;
	wire branchC_59_in1_ready;
	wire branchC_59_in1_valid;
	wire branchC_59_in2_data;
	wire branchC_59_in2_ready;
	wire branchC_59_in2_valid;
	wire branchC_59_out1_data;
	wire branchC_59_out1_ready;
	wire branchC_59_out1_valid;
	wire branchC_59_out2_data;
	wire branchC_59_out2_ready;
	wire branchC_59_out2_valid;
	wire phiC_41_clk;
	wire phiC_41_rst;
	wire phiC_41_in1_data;
	wire phiC_41_in1_ready;
	wire phiC_41_in1_valid;
	wire phiC_41_out1_data;
	wire phiC_41_out1_ready;
	wire phiC_41_out1_valid;
	wire sink_0_clk;
	wire sink_0_rst;
	wire sink_0_in1_data;
	wire sink_0_in1_ready;
	wire sink_0_in1_valid;
	wire sink_1_clk;
	wire sink_1_rst;
	wire [31 : 0] sink_1_in1_data;
	wire sink_1_in1_ready;
	wire sink_1_in1_valid;
	wire sink_2_clk;
	wire sink_2_rst;
	wire [31 : 0] sink_2_in1_data;
	wire sink_2_in1_ready;
	wire sink_2_in1_valid;
	wire sink_3_clk;
	wire sink_3_rst;
	wire sink_3_in1_data;
	wire sink_3_in1_ready;
	wire sink_3_in1_valid;
	wire sink_4_clk;
	wire sink_4_rst;
	wire [5 : 0] sink_4_in1_data;
	wire sink_4_in1_ready;
	wire sink_4_in1_valid;
	wire sink_5_clk;
	wire sink_5_rst;
	wire [31 : 0] sink_5_in1_data;
	wire sink_5_in1_ready;
	wire sink_5_in1_valid;
	wire sink_6_clk;
	wire sink_6_rst;
	wire [31 : 0] sink_6_in1_data;
	wire sink_6_in1_ready;
	wire sink_6_in1_valid;
	wire sink_7_clk;
	wire sink_7_rst;
	wire [5 : 0] sink_7_in1_data;
	wire sink_7_in1_ready;
	wire sink_7_in1_valid;
	wire sink_8_clk;
	wire sink_8_rst;
	wire [5 : 0] sink_8_in1_data;
	wire sink_8_in1_ready;
	wire sink_8_in1_valid;
	wire sink_9_clk;
	wire sink_9_rst;
	wire sink_9_in1_data;
	wire sink_9_in1_ready;
	wire sink_9_in1_valid;
	wire sink_10_clk;
	wire sink_10_rst;
	wire [31 : 0] sink_10_in1_data;
	wire sink_10_in1_ready;
	wire sink_10_in1_valid;
	wire sink_11_clk;
	wire sink_11_rst;
	wire [31 : 0] sink_11_in1_data;
	wire sink_11_in1_ready;
	wire sink_11_in1_valid;
	wire sink_12_clk;
	wire sink_12_rst;
	wire [31 : 0] sink_12_in1_data;
	wire sink_12_in1_ready;
	wire sink_12_in1_valid;
	wire sink_13_clk;
	wire sink_13_rst;
	wire sink_13_in1_data;
	wire sink_13_in1_ready;
	wire sink_13_in1_valid;
	wire sink_14_clk;
	wire sink_14_rst;
	wire [31 : 0] sink_14_in1_data;
	wire sink_14_in1_ready;
	wire sink_14_in1_valid;
	wire sink_15_clk;
	wire sink_15_rst;
	wire [31 : 0] sink_15_in1_data;
	wire sink_15_in1_ready;
	wire sink_15_in1_valid;
	wire sink_16_clk;
	wire sink_16_rst;
	wire [5 : 0] sink_16_in1_data;
	wire sink_16_in1_ready;
	wire sink_16_in1_valid;
	wire sink_17_clk;
	wire sink_17_rst;
	wire [5 : 0] sink_17_in1_data;
	wire sink_17_in1_ready;
	wire sink_17_in1_valid;
	wire sink_18_clk;
	wire sink_18_rst;
	wire [31 : 0] sink_18_in1_data;
	wire sink_18_in1_ready;
	wire sink_18_in1_valid;
	wire sink_19_clk;
	wire sink_19_rst;
	wire [5 : 0] sink_19_in1_data;
	wire sink_19_in1_ready;
	wire sink_19_in1_valid;
	wire sink_20_clk;
	wire sink_20_rst;
	wire sink_20_in1_data;
	wire sink_20_in1_ready;
	wire sink_20_in1_valid;
	wire sink_21_clk;
	wire sink_21_rst;
	wire [31 : 0] sink_21_in1_data;
	wire sink_21_in1_ready;
	wire sink_21_in1_valid;
	wire sink_22_clk;
	wire sink_22_rst;
	wire [5 : 0] sink_22_in1_data;
	wire sink_22_in1_ready;
	wire sink_22_in1_valid;
	wire sink_23_clk;
	wire sink_23_rst;
	wire sink_23_in1_data;
	wire sink_23_in1_ready;
	wire sink_23_in1_valid;
	wire sink_24_clk;
	wire sink_24_rst;
	wire [31 : 0] sink_24_in1_data;
	wire sink_24_in1_ready;
	wire sink_24_in1_valid;
	wire sink_25_clk;
	wire sink_25_rst;
	wire [31 : 0] sink_25_in1_data;
	wire sink_25_in1_ready;
	wire sink_25_in1_valid;
	wire sink_26_clk;
	wire sink_26_rst;
	wire sink_26_in1_data;
	wire sink_26_in1_ready;
	wire sink_26_in1_valid;
	wire sink_27_clk;
	wire sink_27_rst;
	wire [31 : 0] sink_27_in1_data;
	wire sink_27_in1_ready;
	wire sink_27_in1_valid;
	wire sink_28_clk;
	wire sink_28_rst;
	wire [5 : 0] sink_28_in1_data;
	wire sink_28_in1_ready;
	wire sink_28_in1_valid;
	wire sink_29_clk;
	wire sink_29_rst;
	wire [5 : 0] sink_29_in1_data;
	wire sink_29_in1_ready;
	wire sink_29_in1_valid;
	wire sink_30_clk;
	wire sink_30_rst;
	wire [31 : 0] sink_30_in1_data;
	wire sink_30_in1_ready;
	wire sink_30_in1_valid;
	wire sink_31_clk;
	wire sink_31_rst;
	wire [5 : 0] sink_31_in1_data;
	wire sink_31_in1_ready;
	wire sink_31_in1_valid;
	wire sink_32_clk;
	wire sink_32_rst;
	wire sink_32_in1_data;
	wire sink_32_in1_ready;
	wire sink_32_in1_valid;
	wire sink_33_clk;
	wire sink_33_rst;
	wire sink_33_in1_data;
	wire sink_33_in1_ready;
	wire sink_33_in1_valid;
	wire sink_34_clk;
	wire sink_34_rst;
	wire sink_34_in1_data;
	wire sink_34_in1_ready;
	wire sink_34_in1_valid;
	wire sink_35_clk;
	wire sink_35_rst;
	wire sink_35_in1_data;
	wire sink_35_in1_ready;
	wire sink_35_in1_valid;
	wire sink_36_clk;
	wire sink_36_rst;
	wire sink_36_in1_data;
	wire sink_36_in1_ready;
	wire sink_36_in1_valid;
	wire sink_37_clk;
	wire sink_37_rst;
	wire sink_37_in1_data;
	wire sink_37_in1_ready;
	wire sink_37_in1_valid;
	wire sink_38_clk;
	wire sink_38_rst;
	wire sink_38_in1_data;
	wire sink_38_in1_ready;
	wire sink_38_in1_valid;
	wire source_0_clk;
	wire source_0_rst;
	wire [2 : 0] source_0_out1_data;
	wire source_0_out1_ready;
	wire source_0_out1_valid;
	wire source_1_clk;
	wire source_1_rst;
	wire [2 : 0] source_1_out1_data;
	wire source_1_out1_ready;
	wire source_1_out1_valid;
	wire source_2_clk;
	wire source_2_rst;
	wire source_2_out1_data;
	wire source_2_out1_ready;
	wire source_2_out1_valid;
	wire source_3_clk;
	wire source_3_rst;
	wire [5 : 0] source_3_out1_data;
	wire source_3_out1_ready;
	wire source_3_out1_valid;
	wire source_4_clk;
	wire source_4_rst;
	wire source_4_out1_data;
	wire source_4_out1_ready;
	wire source_4_out1_valid;
	wire source_5_clk;
	wire source_5_rst;
	wire [5 : 0] source_5_out1_data;
	wire source_5_out1_ready;
	wire source_5_out1_valid;
	wire source_6_clk;
	wire source_6_rst;
	wire [2 : 0] source_6_out1_data;
	wire source_6_out1_ready;
	wire source_6_out1_valid;
	wire source_7_clk;
	wire source_7_rst;
	wire source_7_out1_data;
	wire source_7_out1_ready;
	wire source_7_out1_valid;
	wire source_8_clk;
	wire source_8_rst;
	wire [5 : 0] source_8_out1_data;
	wire source_8_out1_ready;
	wire source_8_out1_valid;
	wire source_9_clk;
	wire source_9_rst;
	wire source_9_out1_data;
	wire source_9_out1_ready;
	wire source_9_out1_valid;
	wire source_10_clk;
	wire source_10_rst;
	wire [5 : 0] source_10_out1_data;
	wire source_10_out1_ready;
	wire source_10_out1_valid;
	wire source_11_clk;
	wire source_11_rst;
	wire source_11_out1_data;
	wire source_11_out1_ready;
	wire source_11_out1_valid;
	wire source_12_clk;
	wire source_12_rst;
	wire [5 : 0] source_12_out1_data;
	wire source_12_out1_ready;
	wire source_12_out1_valid;
	wire source_13_clk;
	wire source_13_rst;
	wire [2 : 0] source_13_out1_data;
	wire source_13_out1_ready;
	wire source_13_out1_valid;
	wire source_14_clk;
	wire source_14_rst;
	wire source_14_out1_data;
	wire source_14_out1_ready;
	wire source_14_out1_valid;
	wire source_15_clk;
	wire source_15_rst;
	wire [5 : 0] source_15_out1_data;
	wire source_15_out1_ready;
	wire source_15_out1_valid;
	wire source_16_clk;
	wire source_16_rst;
	wire source_16_out1_data;
	wire source_16_out1_ready;
	wire source_16_out1_valid;
	wire source_17_clk;
	wire source_17_rst;
	wire [5 : 0] source_17_out1_data;
	wire source_17_out1_ready;
	wire source_17_out1_valid;
	wire fork_62_clk;
	wire fork_62_rst;
	wire fork_62_in1_data;
	wire fork_62_in1_ready;
	wire fork_62_in1_valid;
	wire fork_62_out1_data;
	wire fork_62_out1_ready;
	wire fork_62_out1_valid;
	wire fork_62_out2_data;
	wire fork_62_out2_ready;
	wire fork_62_out2_valid;
	wire fork_65_clk;
	wire fork_65_rst;
	wire fork_65_in1_data;
	wire fork_65_in1_ready;
	wire fork_65_in1_valid;
	wire fork_65_out1_data;
	wire fork_65_out1_ready;
	wire fork_65_out1_valid;
	wire fork_65_out2_data;
	wire fork_65_out2_ready;
	wire fork_65_out2_valid;
	wire Buffer_0_clk;
	wire Buffer_0_rst;
	wire [5 : 0] Buffer_0_in1_data;
	wire Buffer_0_in1_ready;
	wire Buffer_0_in1_valid;
	wire [5 : 0] Buffer_0_out1_data;
	wire Buffer_0_out1_ready;
	wire Buffer_0_out1_valid;
	wire Buffer_1_clk;
	wire Buffer_1_rst;
	wire [31 : 0] Buffer_1_in1_data;
	wire Buffer_1_in1_ready;
	wire Buffer_1_in1_valid;
	wire [31 : 0] Buffer_1_out1_data;
	wire Buffer_1_out1_ready;
	wire Buffer_1_out1_valid;
	wire Buffer_2_clk;
	wire Buffer_2_rst;
	wire Buffer_2_in1_data;
	wire Buffer_2_in1_ready;
	wire Buffer_2_in1_valid;
	wire Buffer_2_out1_data;
	wire Buffer_2_out1_ready;
	wire Buffer_2_out1_valid;
	wire Buffer_3_clk;
	wire Buffer_3_rst;
	wire [5 : 0] Buffer_3_in1_data;
	wire Buffer_3_in1_ready;
	wire Buffer_3_in1_valid;
	wire [5 : 0] Buffer_3_out1_data;
	wire Buffer_3_out1_ready;
	wire Buffer_3_out1_valid;
	wire Buffer_4_clk;
	wire Buffer_4_rst;
	wire [31 : 0] Buffer_4_in1_data;
	wire Buffer_4_in1_ready;
	wire Buffer_4_in1_valid;
	wire [31 : 0] Buffer_4_out1_data;
	wire Buffer_4_out1_ready;
	wire Buffer_4_out1_valid;
	wire Buffer_5_clk;
	wire Buffer_5_rst;
	wire [31 : 0] Buffer_5_in1_data;
	wire Buffer_5_in1_ready;
	wire Buffer_5_in1_valid;
	wire [31 : 0] Buffer_5_out1_data;
	wire Buffer_5_out1_ready;
	wire Buffer_5_out1_valid;
	wire Buffer_6_clk;
	wire Buffer_6_rst;
	wire Buffer_6_in1_data;
	wire Buffer_6_in1_ready;
	wire Buffer_6_in1_valid;
	wire Buffer_6_out1_data;
	wire Buffer_6_out1_ready;
	wire Buffer_6_out1_valid;
	wire Buffer_7_clk;
	wire Buffer_7_rst;
	wire Buffer_7_in1_data;
	wire Buffer_7_in1_ready;
	wire Buffer_7_in1_valid;
	wire Buffer_7_out1_data;
	wire Buffer_7_out1_ready;
	wire Buffer_7_out1_valid;
	wire Buffer_8_clk;
	wire Buffer_8_rst;
	wire [31 : 0] Buffer_8_in1_data;
	wire Buffer_8_in1_ready;
	wire Buffer_8_in1_valid;
	wire [31 : 0] Buffer_8_out1_data;
	wire Buffer_8_out1_ready;
	wire Buffer_8_out1_valid;
	wire Buffer_9_clk;
	wire Buffer_9_rst;
	wire [5 : 0] Buffer_9_in1_data;
	wire Buffer_9_in1_ready;
	wire Buffer_9_in1_valid;
	wire [5 : 0] Buffer_9_out1_data;
	wire Buffer_9_out1_ready;
	wire Buffer_9_out1_valid;
	wire Buffer_10_clk;
	wire Buffer_10_rst;
	wire [5 : 0] Buffer_10_in1_data;
	wire Buffer_10_in1_ready;
	wire Buffer_10_in1_valid;
	wire [5 : 0] Buffer_10_out1_data;
	wire Buffer_10_out1_ready;
	wire Buffer_10_out1_valid;
	wire Buffer_11_clk;
	wire Buffer_11_rst;
	wire [31 : 0] Buffer_11_in1_data;
	wire Buffer_11_in1_ready;
	wire Buffer_11_in1_valid;
	wire [31 : 0] Buffer_11_out1_data;
	wire Buffer_11_out1_ready;
	wire Buffer_11_out1_valid;
	wire Buffer_12_clk;
	wire Buffer_12_rst;
	wire [31 : 0] Buffer_12_in1_data;
	wire Buffer_12_in1_ready;
	wire Buffer_12_in1_valid;
	wire [31 : 0] Buffer_12_out1_data;
	wire Buffer_12_out1_ready;
	wire Buffer_12_out1_valid;
	wire Buffer_13_clk;
	wire Buffer_13_rst;
	wire [31 : 0] Buffer_13_in1_data;
	wire Buffer_13_in1_ready;
	wire Buffer_13_in1_valid;
	wire [31 : 0] Buffer_13_out1_data;
	wire Buffer_13_out1_ready;
	wire Buffer_13_out1_valid;
	wire Buffer_14_clk;
	wire Buffer_14_rst;
	wire [5 : 0] Buffer_14_in1_data;
	wire Buffer_14_in1_ready;
	wire Buffer_14_in1_valid;
	wire [5 : 0] Buffer_14_out1_data;
	wire Buffer_14_out1_ready;
	wire Buffer_14_out1_valid;
	wire Buffer_15_clk;
	wire Buffer_15_rst;
	wire [5 : 0] Buffer_15_in1_data;
	wire Buffer_15_in1_ready;
	wire Buffer_15_in1_valid;
	wire [5 : 0] Buffer_15_out1_data;
	wire Buffer_15_out1_ready;
	wire Buffer_15_out1_valid;
	wire Buffer_16_clk;
	wire Buffer_16_rst;
	wire Buffer_16_in1_data;
	wire Buffer_16_in1_ready;
	wire Buffer_16_in1_valid;
	wire Buffer_16_out1_data;
	wire Buffer_16_out1_ready;
	wire Buffer_16_out1_valid;
	wire Buffer_17_clk;
	wire Buffer_17_rst;
	wire [5 : 0] Buffer_17_in1_data;
	wire Buffer_17_in1_ready;
	wire Buffer_17_in1_valid;
	wire [5 : 0] Buffer_17_out1_data;
	wire Buffer_17_out1_ready;
	wire Buffer_17_out1_valid;
	wire Buffer_18_clk;
	wire Buffer_18_rst;
	wire [31 : 0] Buffer_18_in1_data;
	wire Buffer_18_in1_ready;
	wire Buffer_18_in1_valid;
	wire [31 : 0] Buffer_18_out1_data;
	wire Buffer_18_out1_ready;
	wire Buffer_18_out1_valid;
	wire Buffer_19_clk;
	wire Buffer_19_rst;
	wire [31 : 0] Buffer_19_in1_data;
	wire Buffer_19_in1_ready;
	wire Buffer_19_in1_valid;
	wire [31 : 0] Buffer_19_out1_data;
	wire Buffer_19_out1_ready;
	wire Buffer_19_out1_valid;
	wire Buffer_20_clk;
	wire Buffer_20_rst;
	wire Buffer_20_in1_data;
	wire Buffer_20_in1_ready;
	wire Buffer_20_in1_valid;
	wire Buffer_20_out1_data;
	wire Buffer_20_out1_ready;
	wire Buffer_20_out1_valid;
	wire Buffer_21_clk;
	wire Buffer_21_rst;
	wire Buffer_21_in1_data;
	wire Buffer_21_in1_ready;
	wire Buffer_21_in1_valid;
	wire Buffer_21_out1_data;
	wire Buffer_21_out1_ready;
	wire Buffer_21_out1_valid;
	wire Buffer_22_clk;
	wire Buffer_22_rst;
	wire [31 : 0] Buffer_22_in1_data;
	wire Buffer_22_in1_ready;
	wire Buffer_22_in1_valid;
	wire [31 : 0] Buffer_22_out1_data;
	wire Buffer_22_out1_ready;
	wire Buffer_22_out1_valid;
	wire Buffer_23_clk;
	wire Buffer_23_rst;
	wire [31 : 0] Buffer_23_in1_data;
	wire Buffer_23_in1_ready;
	wire Buffer_23_in1_valid;
	wire [31 : 0] Buffer_23_out1_data;
	wire Buffer_23_out1_ready;
	wire Buffer_23_out1_valid;
	wire Buffer_24_clk;
	wire Buffer_24_rst;
	wire [31 : 0] Buffer_24_in1_data;
	wire Buffer_24_in1_ready;
	wire Buffer_24_in1_valid;
	wire [31 : 0] Buffer_24_out1_data;
	wire Buffer_24_out1_ready;
	wire Buffer_24_out1_valid;
	wire Buffer_25_clk;
	wire Buffer_25_rst;
	wire [5 : 0] Buffer_25_in1_data;
	wire Buffer_25_in1_ready;
	wire Buffer_25_in1_valid;
	wire [5 : 0] Buffer_25_out1_data;
	wire Buffer_25_out1_ready;
	wire Buffer_25_out1_valid;
	wire Buffer_26_clk;
	wire Buffer_26_rst;
	wire [5 : 0] Buffer_26_in1_data;
	wire Buffer_26_in1_ready;
	wire Buffer_26_in1_valid;
	wire [5 : 0] Buffer_26_out1_data;
	wire Buffer_26_out1_ready;
	wire Buffer_26_out1_valid;
	wire Buffer_27_clk;
	wire Buffer_27_rst;
	wire Buffer_27_in1_data;
	wire Buffer_27_in1_ready;
	wire Buffer_27_in1_valid;
	wire Buffer_27_out1_data;
	wire Buffer_27_out1_ready;
	wire Buffer_27_out1_valid;
	wire Buffer_28_clk;
	wire Buffer_28_rst;
	wire [31 : 0] Buffer_28_in1_data;
	wire Buffer_28_in1_ready;
	wire Buffer_28_in1_valid;
	wire [31 : 0] Buffer_28_out1_data;
	wire Buffer_28_out1_ready;
	wire Buffer_28_out1_valid;
	wire Buffer_29_clk;
	wire Buffer_29_rst;
	wire [5 : 0] Buffer_29_in1_data;
	wire Buffer_29_in1_ready;
	wire Buffer_29_in1_valid;
	wire [5 : 0] Buffer_29_out1_data;
	wire Buffer_29_out1_ready;
	wire Buffer_29_out1_valid;
	assign Buffer_30_clk = clk;
	assign Buffer_30_rst = rst;
	assign forkC_55_in1_data = Buffer_30__forkC_55__data__0__anchor__in;
	assign Buffer_30__forkC_55__data__0__anchor__out = Buffer_30_out1_data;
	assign forkC_55_in1_valid = Buffer_30__forkC_55__valid__0__anchor__in;
	assign Buffer_30__forkC_55__valid__0__anchor__out = Buffer_30_out1_valid;
	assign Buffer_30_out1_ready = Buffer_30__forkC_55__ready__0__anchor__in;
	assign Buffer_30__forkC_55__ready__0__anchor__out = forkC_55_in1_ready;
	assign alpha_clk = clk;
	assign alpha_rst = rst;
	assign alpha_in1_data = alpha_din;
	assign alpha_in1_valid = alpha_valid_in;
	assign alpha_ready_in = alpha_in1_ready;
	assign branch_2_in1_data = alpha__branch_2__data__0__anchor__in;
	assign alpha__branch_2__data__0__anchor__out = alpha_out1_data;
	assign branch_2_in1_valid = alpha__branch_2__valid__0__anchor__in;
	assign alpha__branch_2__valid__0__anchor__out = alpha_out1_valid;
	assign alpha_out1_ready = alpha__branch_2__ready__0__anchor__in;
	assign alpha__branch_2__ready__0__anchor__out = branch_2_in1_ready;
	assign beta_clk = clk;
	assign beta_rst = rst;
	assign beta_in1_data = beta_din;
	assign beta_in1_valid = beta_valid_in;
	assign beta_ready_in = beta_in1_ready;
	assign branch_1_in1_data = beta__branch_1__data__0__anchor__in;
	assign beta__branch_1__data__0__anchor__out = beta_out1_data;
	assign branch_1_in1_valid = beta__branch_1__valid__0__anchor__in;
	assign beta__branch_1__valid__0__anchor__out = beta_out1_valid;
	assign beta_out1_ready = beta__branch_1__ready__0__anchor__in;
	assign beta__branch_1__ready__0__anchor__out = branch_1_in1_ready;
	assign brCst_block1_clk = clk;
	assign brCst_block1_rst = rst;
	assign fork_29_in1_data = brCst_block1__fork_29__data__0__anchor__in;
	assign brCst_block1__fork_29__data__0__anchor__out = brCst_block1_out1_data;
	assign fork_29_in1_valid = brCst_block1__fork_29__valid__0__anchor__in;
	assign brCst_block1__fork_29__valid__0__anchor__out = brCst_block1_out1_valid;
	assign brCst_block1_out1_ready = brCst_block1__fork_29__ready__0__anchor__in;
	assign brCst_block1__fork_29__ready__0__anchor__out = fork_29_in1_ready;
	assign cst_0_clk = clk;
	assign cst_0_rst = rst;
	assign branch_0_in1_data = cst_0__branch_0__data__0__anchor__in;
	assign cst_0__branch_0__data__0__anchor__out = cst_0_out1_data;
	assign branch_0_in1_valid = cst_0__branch_0__valid__0__anchor__in;
	assign cst_0__branch_0__valid__0__anchor__out = cst_0_out1_valid;
	assign cst_0_out1_ready = cst_0__branch_0__ready__0__anchor__in;
	assign cst_0__branch_0__ready__0__anchor__out = branch_0_in1_ready;
	assign phi_1_clk = clk;
	assign phi_1_rst = rst;
	assign branch_4_in1_data = phi_1__branch_4__data__0__anchor__in;
	assign phi_1__branch_4__data__0__anchor__out = phi_1_out1_data;
	assign branch_4_in1_valid = phi_1__branch_4__valid__0__anchor__in;
	assign phi_1__branch_4__valid__0__anchor__out = phi_1_out1_valid;
	assign phi_1_out1_ready = phi_1__branch_4__ready__0__anchor__in;
	assign phi_1__branch_4__ready__0__anchor__out = branch_4_in1_ready;
	assign brCst_block2_clk = clk;
	assign brCst_block2_rst = rst;
	assign fork_30_in1_data = brCst_block2__fork_30__data__0__anchor__in;
	assign brCst_block2__fork_30__data__0__anchor__out = brCst_block2_out1_data;
	assign fork_30_in1_valid = brCst_block2__fork_30__valid__0__anchor__in;
	assign brCst_block2__fork_30__valid__0__anchor__out = brCst_block2_out1_valid;
	assign brCst_block2_out1_ready = brCst_block2__fork_30__ready__0__anchor__in;
	assign brCst_block2__fork_30__ready__0__anchor__out = fork_30_in1_ready;
	assign cst_1_clk = clk;
	assign cst_1_rst = rst;
	assign branch_3_in1_data = cst_1__branch_3__data__0__anchor__in;
	assign cst_1__branch_3__data__0__anchor__out = cst_1_out1_data;
	assign branch_3_in1_valid = cst_1__branch_3__valid__0__anchor__in;
	assign cst_1__branch_3__valid__0__anchor__out = cst_1_out1_valid;
	assign cst_1_out1_ready = cst_1__branch_3__ready__0__anchor__in;
	assign cst_1__branch_3__ready__0__anchor__out = branch_3_in1_ready;
	assign phi_3_clk = clk;
	assign phi_3_rst = rst;
	assign fork_0_in1_data = phi_3__fork_0__data__0__anchor__in;
	assign phi_3__fork_0__data__0__anchor__out = phi_3_out1_data;
	assign fork_0_in1_valid = phi_3__fork_0__valid__0__anchor__in;
	assign phi_3__fork_0__valid__0__anchor__out = phi_3_out1_valid;
	assign phi_3_out1_ready = phi_3__fork_0__ready__0__anchor__in;
	assign phi_3__fork_0__ready__0__anchor__out = fork_0_in1_ready;
	assign cst_2_clk = clk;
	assign cst_2_rst = rst;
	assign shl_4_in2_data = cst_2__shl_4__data__0__anchor__in;
	assign cst_2__shl_4__data__0__anchor__out = cst_2_out1_data;
	assign shl_4_in2_valid = cst_2__shl_4__valid__0__anchor__in;
	assign cst_2__shl_4__valid__0__anchor__out = cst_2_out1_valid;
	assign cst_2_out1_ready = cst_2__shl_4__ready__0__anchor__in;
	assign cst_2__shl_4__ready__0__anchor__out = shl_4_in2_ready;
	assign shl_4_clk = clk;
	assign shl_4_rst = rst;
	assign add_5_in1_data = shl_4__add_5__data__0__anchor__in;
	assign shl_4__add_5__data__0__anchor__out = shl_4_out1_data;
	assign add_5_in1_valid = shl_4__add_5__valid__0__anchor__in;
	assign shl_4__add_5__valid__0__anchor__out = shl_4_out1_valid;
	assign shl_4_out1_ready = shl_4__add_5__ready__0__anchor__in;
	assign shl_4__add_5__ready__0__anchor__out = add_5_in1_ready;
	assign add_5_clk = clk;
	assign add_5_rst = rst;
	assign load_8_in2_data = add_5__load_8__data__0__anchor__in;
	assign add_5__load_8__data__0__anchor__out = add_5_out1_data;
	assign load_8_in2_valid = add_5__load_8__valid__0__anchor__in;
	assign add_5__load_8__valid__0__anchor__out = add_5_out1_valid;
	assign add_5_out1_ready = add_5__load_8__ready__0__anchor__in;
	assign add_5__load_8__ready__0__anchor__out = load_8_in2_ready;
	assign load_8_clk = clk;
	assign load_8_rst = rst;
	assign add_16_in1_data = load_8__add_16__data__0__anchor__in;
	assign load_8__add_16__data__0__anchor__out = load_8_out1_data;
	assign add_16_in1_valid = load_8__add_16__valid__0__anchor__in;
	assign load_8__add_16__valid__0__anchor__out = load_8_out1_valid;
	assign load_8_out1_ready = load_8__add_16__ready__0__anchor__in;
	assign load_8__add_16__ready__0__anchor__out = add_16_in1_ready;
	assign MC_A_in2_data = load_8__MC_A__data__0__anchor__in;
	assign load_8__MC_A__data__0__anchor__out = load_8_out2_data;
	assign MC_A_in2_valid = load_8__MC_A__valid__0__anchor__in;
	assign load_8__MC_A__valid__0__anchor__out = load_8_out2_valid;
	assign load_8_out2_ready = load_8__MC_A__ready__0__anchor__in;
	assign load_8__MC_A__ready__0__anchor__out = MC_A_in2_ready;
	assign load_11_clk = clk;
	assign load_11_rst = rst;
	assign mul_15_in1_data = load_11__mul_15__data__0__anchor__in;
	assign load_11__mul_15__data__0__anchor__out = load_11_out1_data;
	assign mul_15_in1_valid = load_11__mul_15__valid__0__anchor__in;
	assign load_11__mul_15__valid__0__anchor__out = load_11_out1_valid;
	assign load_11_out1_ready = load_11__mul_15__ready__0__anchor__in;
	assign load_11__mul_15__ready__0__anchor__out = mul_15_in1_ready;
	assign MC_u1_in1_data = load_11__MC_u1__data__0__anchor__in;
	assign load_11__MC_u1__data__0__anchor__out = load_11_out2_data;
	assign MC_u1_in1_valid = load_11__MC_u1__valid__0__anchor__in;
	assign load_11__MC_u1__valid__0__anchor__out = load_11_out2_valid;
	assign load_11_out2_ready = load_11__MC_u1__ready__0__anchor__in;
	assign load_11__MC_u1__ready__0__anchor__out = MC_u1_in1_ready;
	assign load_14_clk = clk;
	assign load_14_rst = rst;
	assign mul_15_in2_data = load_14__mul_15__data__0__anchor__in;
	assign load_14__mul_15__data__0__anchor__out = load_14_out1_data;
	assign mul_15_in2_valid = load_14__mul_15__valid__0__anchor__in;
	assign load_14__mul_15__valid__0__anchor__out = load_14_out1_valid;
	assign load_14_out1_ready = load_14__mul_15__ready__0__anchor__in;
	assign load_14__mul_15__ready__0__anchor__out = mul_15_in2_ready;
	assign MC_v1_in1_data = load_14__MC_v1__data__0__anchor__in;
	assign load_14__MC_v1__data__0__anchor__out = load_14_out2_data;
	assign MC_v1_in1_valid = load_14__MC_v1__valid__0__anchor__in;
	assign load_14__MC_v1__valid__0__anchor__out = load_14_out2_valid;
	assign load_14_out2_ready = load_14__MC_v1__ready__0__anchor__in;
	assign load_14__MC_v1__ready__0__anchor__out = MC_v1_in1_ready;
	assign mul_15_clk = clk;
	assign mul_15_rst = rst;
	assign add_16_in2_data = mul_15__add_16__data__0__anchor__in;
	assign mul_15__add_16__data__0__anchor__out = mul_15_out1_data;
	assign add_16_in2_valid = mul_15__add_16__valid__0__anchor__in;
	assign mul_15__add_16__valid__0__anchor__out = mul_15_out1_valid;
	assign mul_15_out1_ready = mul_15__add_16__ready__0__anchor__in;
	assign mul_15__add_16__ready__0__anchor__out = add_16_in2_ready;
	assign add_16_clk = clk;
	assign add_16_rst = rst;
	assign add_24_in1_data = add_16__add_24__data__0__anchor__in;
	assign add_16__add_24__data__0__anchor__out = add_16_out1_data;
	assign add_24_in1_valid = add_16__add_24__valid__0__anchor__in;
	assign add_16__add_24__valid__0__anchor__out = add_16_out1_valid;
	assign add_16_out1_ready = add_16__add_24__ready__0__anchor__in;
	assign add_16__add_24__ready__0__anchor__out = add_24_in1_ready;
	assign load_19_clk = clk;
	assign load_19_rst = rst;
	assign mul_23_in1_data = load_19__mul_23__data__0__anchor__in;
	assign load_19__mul_23__data__0__anchor__out = load_19_out1_data;
	assign mul_23_in1_valid = load_19__mul_23__valid__0__anchor__in;
	assign load_19__mul_23__valid__0__anchor__out = load_19_out1_valid;
	assign load_19_out1_ready = load_19__mul_23__ready__0__anchor__in;
	assign load_19__mul_23__ready__0__anchor__out = mul_23_in1_ready;
	assign MC_u2_in1_data = load_19__MC_u2__data__0__anchor__in;
	assign load_19__MC_u2__data__0__anchor__out = load_19_out2_data;
	assign MC_u2_in1_valid = load_19__MC_u2__valid__0__anchor__in;
	assign load_19__MC_u2__valid__0__anchor__out = load_19_out2_valid;
	assign load_19_out2_ready = load_19__MC_u2__ready__0__anchor__in;
	assign load_19__MC_u2__ready__0__anchor__out = MC_u2_in1_ready;
	assign load_22_clk = clk;
	assign load_22_rst = rst;
	assign mul_23_in2_data = load_22__mul_23__data__0__anchor__in;
	assign load_22__mul_23__data__0__anchor__out = load_22_out1_data;
	assign mul_23_in2_valid = load_22__mul_23__valid__0__anchor__in;
	assign load_22__mul_23__valid__0__anchor__out = load_22_out1_valid;
	assign load_22_out1_ready = load_22__mul_23__ready__0__anchor__in;
	assign load_22__mul_23__ready__0__anchor__out = mul_23_in2_ready;
	assign MC_v2_in1_data = load_22__MC_v2__data__0__anchor__in;
	assign load_22__MC_v2__data__0__anchor__out = load_22_out2_data;
	assign MC_v2_in1_valid = load_22__MC_v2__valid__0__anchor__in;
	assign load_22__MC_v2__valid__0__anchor__out = load_22_out2_valid;
	assign load_22_out2_ready = load_22__MC_v2__ready__0__anchor__in;
	assign load_22__MC_v2__ready__0__anchor__out = MC_v2_in1_ready;
	assign mul_23_clk = clk;
	assign mul_23_rst = rst;
	assign add_24_in2_data = mul_23__add_24__data__0__anchor__in;
	assign mul_23__add_24__data__0__anchor__out = mul_23_out1_data;
	assign add_24_in2_valid = mul_23__add_24__valid__0__anchor__in;
	assign mul_23__add_24__valid__0__anchor__out = mul_23_out1_valid;
	assign mul_23_out1_ready = mul_23__add_24__ready__0__anchor__in;
	assign mul_23__add_24__ready__0__anchor__out = add_24_in2_ready;
	assign add_24_clk = clk;
	assign add_24_rst = rst;
	assign store_0_in1_data = add_24__store_0__data__0__anchor__in;
	assign add_24__store_0__data__0__anchor__out = add_24_out1_data;
	assign store_0_in1_valid = add_24__store_0__valid__0__anchor__in;
	assign add_24__store_0__valid__0__anchor__out = add_24_out1_valid;
	assign add_24_out1_ready = add_24__store_0__ready__0__anchor__in;
	assign add_24__store_0__ready__0__anchor__out = store_0_in1_ready;
	assign cst_3_clk = clk;
	assign cst_3_rst = rst;
	assign shl_25_in2_data = cst_3__shl_25__data__0__anchor__in;
	assign cst_3__shl_25__data__0__anchor__out = cst_3_out1_data;
	assign shl_25_in2_valid = cst_3__shl_25__valid__0__anchor__in;
	assign cst_3__shl_25__valid__0__anchor__out = cst_3_out1_valid;
	assign cst_3_out1_ready = cst_3__shl_25__ready__0__anchor__in;
	assign cst_3__shl_25__ready__0__anchor__out = shl_25_in2_ready;
	assign shl_25_clk = clk;
	assign shl_25_rst = rst;
	assign add_26_in1_data = shl_25__add_26__data__0__anchor__in;
	assign shl_25__add_26__data__0__anchor__out = shl_25_out1_data;
	assign add_26_in1_valid = shl_25__add_26__valid__0__anchor__in;
	assign shl_25__add_26__valid__0__anchor__out = shl_25_out1_valid;
	assign shl_25_out1_ready = shl_25__add_26__ready__0__anchor__in;
	assign shl_25__add_26__ready__0__anchor__out = add_26_in1_ready;
	assign add_26_clk = clk;
	assign add_26_rst = rst;
	assign store_0_in2_data = add_26__store_0__data__0__anchor__in;
	assign add_26__store_0__data__0__anchor__out = add_26_out1_data;
	assign store_0_in2_valid = add_26__store_0__valid__0__anchor__in;
	assign add_26__store_0__valid__0__anchor__out = add_26_out1_valid;
	assign add_26_out1_ready = add_26__store_0__ready__0__anchor__in;
	assign add_26__store_0__ready__0__anchor__out = store_0_in2_ready;
	assign store_0_clk = clk;
	assign store_0_rst = rst;
	assign MC_A_in4_data = store_0__MC_A__data__0__anchor__in;
	assign store_0__MC_A__data__0__anchor__out = store_0_out1_data;
	assign MC_A_in4_valid = store_0__MC_A__valid__0__anchor__in;
	assign store_0__MC_A__valid__0__anchor__out = store_0_out1_valid;
	assign store_0_out1_ready = store_0__MC_A__ready__0__anchor__in;
	assign store_0__MC_A__ready__0__anchor__out = MC_A_in4_ready;
	assign MC_A_in3_data = store_0__MC_A__data__1__anchor__in;
	assign store_0__MC_A__data__1__anchor__out = store_0_out2_data;
	assign MC_A_in3_valid = store_0__MC_A__valid__1__anchor__in;
	assign store_0__MC_A__valid__1__anchor__out = store_0_out2_valid;
	assign store_0_out2_ready = store_0__MC_A__ready__1__anchor__in;
	assign store_0__MC_A__ready__1__anchor__out = MC_A_in3_ready;
	assign cst_4_clk = clk;
	assign cst_4_rst = rst;
	assign add_29_in2_data = cst_4__add_29__data__0__anchor__in;
	assign cst_4__add_29__data__0__anchor__out = cst_4_out1_data;
	assign add_29_in2_valid = cst_4__add_29__valid__0__anchor__in;
	assign cst_4__add_29__valid__0__anchor__out = cst_4_out1_valid;
	assign cst_4_out1_ready = cst_4__add_29__ready__0__anchor__in;
	assign cst_4__add_29__ready__0__anchor__out = add_29_in2_ready;
	assign add_29_clk = clk;
	assign add_29_rst = rst;
	assign fork_1_in1_data = add_29__fork_1__data__0__anchor__in;
	assign add_29__fork_1__data__0__anchor__out = add_29_out1_data;
	assign fork_1_in1_valid = add_29__fork_1__valid__0__anchor__in;
	assign add_29__fork_1__valid__0__anchor__out = add_29_out1_valid;
	assign add_29_out1_ready = add_29__fork_1__ready__0__anchor__in;
	assign add_29__fork_1__ready__0__anchor__out = fork_1_in1_ready;
	assign cst_5_clk = clk;
	assign cst_5_rst = rst;
	assign icmp_30_in2_data = cst_5__icmp_30__data__0__anchor__in;
	assign cst_5__icmp_30__data__0__anchor__out = cst_5_out1_data;
	assign icmp_30_in2_valid = cst_5__icmp_30__valid__0__anchor__in;
	assign cst_5__icmp_30__valid__0__anchor__out = cst_5_out1_valid;
	assign cst_5_out1_ready = cst_5__icmp_30__ready__0__anchor__in;
	assign cst_5__icmp_30__ready__0__anchor__out = icmp_30_in2_ready;
	assign icmp_30_clk = clk;
	assign icmp_30_rst = rst;
	assign fork_31_in1_data = icmp_30__fork_31__data__0__anchor__in;
	assign icmp_30__fork_31__data__0__anchor__out = icmp_30_out1_data;
	assign fork_31_in1_valid = icmp_30__fork_31__valid__0__anchor__in;
	assign icmp_30__fork_31__valid__0__anchor__out = icmp_30_out1_valid;
	assign icmp_30_out1_ready = icmp_30__fork_31__ready__0__anchor__in;
	assign icmp_30__fork_31__ready__0__anchor__out = fork_31_in1_ready;
	assign cst_6_clk = clk;
	assign cst_6_rst = rst;
	assign add_32_in2_data = cst_6__add_32__data__0__anchor__in;
	assign cst_6__add_32__data__0__anchor__out = cst_6_out1_data;
	assign add_32_in2_valid = cst_6__add_32__valid__0__anchor__in;
	assign cst_6__add_32__valid__0__anchor__out = cst_6_out1_valid;
	assign cst_6_out1_ready = cst_6__add_32__ready__0__anchor__in;
	assign cst_6__add_32__ready__0__anchor__out = add_32_in2_ready;
	assign add_32_clk = clk;
	assign add_32_rst = rst;
	assign fork_2_in1_data = add_32__fork_2__data__0__anchor__in;
	assign add_32__fork_2__data__0__anchor__out = add_32_out1_data;
	assign fork_2_in1_valid = add_32__fork_2__valid__0__anchor__in;
	assign add_32__fork_2__valid__0__anchor__out = add_32_out1_valid;
	assign add_32_out1_ready = add_32__fork_2__ready__0__anchor__in;
	assign add_32__fork_2__ready__0__anchor__out = fork_2_in1_ready;
	assign cst_7_clk = clk;
	assign cst_7_rst = rst;
	assign icmp_33_in2_data = cst_7__icmp_33__data__0__anchor__in;
	assign cst_7__icmp_33__data__0__anchor__out = cst_7_out1_data;
	assign icmp_33_in2_valid = cst_7__icmp_33__valid__0__anchor__in;
	assign cst_7__icmp_33__valid__0__anchor__out = cst_7_out1_valid;
	assign cst_7_out1_ready = cst_7__icmp_33__ready__0__anchor__in;
	assign cst_7__icmp_33__ready__0__anchor__out = icmp_33_in2_ready;
	assign icmp_33_clk = clk;
	assign icmp_33_rst = rst;
	assign fork_32_in1_data = icmp_33__fork_32__data__0__anchor__in;
	assign icmp_33__fork_32__data__0__anchor__out = icmp_33_out1_data;
	assign fork_32_in1_valid = icmp_33__fork_32__valid__0__anchor__in;
	assign icmp_33__fork_32__valid__0__anchor__out = icmp_33_out1_valid;
	assign icmp_33_out1_ready = icmp_33__fork_32__ready__0__anchor__in;
	assign icmp_33__fork_32__ready__0__anchor__out = fork_32_in1_ready;
	assign brCst_block5_clk = clk;
	assign brCst_block5_rst = rst;
	assign fork_33_in1_data = brCst_block5__fork_33__data__0__anchor__in;
	assign brCst_block5__fork_33__data__0__anchor__out = brCst_block5_out1_data;
	assign fork_33_in1_valid = brCst_block5__fork_33__valid__0__anchor__in;
	assign brCst_block5__fork_33__valid__0__anchor__out = brCst_block5_out1_valid;
	assign brCst_block5_out1_ready = brCst_block5__fork_33__ready__0__anchor__in;
	assign brCst_block5__fork_33__ready__0__anchor__out = fork_33_in1_ready;
	assign cst_8_clk = clk;
	assign cst_8_rst = rst;
	assign branch_14_in1_data = cst_8__branch_14__data__0__anchor__in;
	assign cst_8__branch_14__data__0__anchor__out = cst_8_out1_data;
	assign branch_14_in1_valid = cst_8__branch_14__valid__0__anchor__in;
	assign cst_8__branch_14__valid__0__anchor__out = cst_8_out1_valid;
	assign cst_8_out1_ready = cst_8__branch_14__ready__0__anchor__in;
	assign cst_8__branch_14__ready__0__anchor__out = branch_14_in1_ready;
	assign phi_36_clk = clk;
	assign phi_36_rst = rst;
	assign fork_3_in1_data = phi_36__fork_3__data__0__anchor__in;
	assign phi_36__fork_3__data__0__anchor__out = phi_36_out1_data;
	assign fork_3_in1_valid = phi_36__fork_3__valid__0__anchor__in;
	assign phi_36__fork_3__valid__0__anchor__out = phi_36_out1_valid;
	assign phi_36_out1_ready = phi_36__fork_3__ready__0__anchor__in;
	assign phi_36__fork_3__ready__0__anchor__out = fork_3_in1_ready;
	assign load_39_clk = clk;
	assign load_39_rst = rst;
	assign branch_17_in1_data = load_39__branch_17__data__0__anchor__in;
	assign load_39__branch_17__data__0__anchor__out = load_39_out1_data;
	assign branch_17_in1_valid = load_39__branch_17__valid__0__anchor__in;
	assign load_39__branch_17__valid__0__anchor__out = load_39_out1_valid;
	assign load_39_out1_ready = load_39__branch_17__ready__0__anchor__in;
	assign load_39__branch_17__ready__0__anchor__out = branch_17_in1_ready;
	assign MC_x_in3_data = load_39__MC_x__data__0__anchor__in;
	assign load_39__MC_x__data__0__anchor__out = load_39_out2_data;
	assign MC_x_in3_valid = load_39__MC_x__valid__0__anchor__in;
	assign load_39__MC_x__valid__0__anchor__out = load_39_out2_valid;
	assign load_39_out2_ready = load_39__MC_x__ready__0__anchor__in;
	assign load_39__MC_x__ready__0__anchor__out = MC_x_in3_ready;
	assign brCst_block6_clk = clk;
	assign brCst_block6_rst = rst;
	assign fork_34_in1_data = brCst_block6__fork_34__data__0__anchor__in;
	assign brCst_block6__fork_34__data__0__anchor__out = brCst_block6_out1_data;
	assign fork_34_in1_valid = brCst_block6__fork_34__valid__0__anchor__in;
	assign brCst_block6__fork_34__valid__0__anchor__out = brCst_block6_out1_valid;
	assign brCst_block6_out1_ready = brCst_block6__fork_34__ready__0__anchor__in;
	assign brCst_block6__fork_34__ready__0__anchor__out = fork_34_in1_ready;
	assign phi_41_clk = clk;
	assign phi_41_rst = rst;
	assign add_53_in1_data = phi_41__add_53__data__0__anchor__in;
	assign phi_41__add_53__data__0__anchor__out = phi_41_out1_data;
	assign add_53_in1_valid = phi_41__add_53__valid__0__anchor__in;
	assign phi_41__add_53__valid__0__anchor__out = phi_41_out1_valid;
	assign phi_41_out1_ready = phi_41__add_53__ready__0__anchor__in;
	assign phi_41__add_53__ready__0__anchor__out = add_53_in1_ready;
	assign cst_9_clk = clk;
	assign cst_9_rst = rst;
	assign branch_18_in1_data = cst_9__branch_18__data__0__anchor__in;
	assign cst_9__branch_18__data__0__anchor__out = cst_9_out1_data;
	assign branch_18_in1_valid = cst_9__branch_18__valid__0__anchor__in;
	assign cst_9__branch_18__valid__0__anchor__out = cst_9_out1_valid;
	assign cst_9_out1_ready = cst_9__branch_18__ready__0__anchor__in;
	assign cst_9__branch_18__ready__0__anchor__out = branch_18_in1_ready;
	assign phi_42_clk = clk;
	assign phi_42_rst = rst;
	assign fork_4_in1_data = phi_42__fork_4__data__0__anchor__in;
	assign phi_42__fork_4__data__0__anchor__out = phi_42_out1_data;
	assign fork_4_in1_valid = phi_42__fork_4__valid__0__anchor__in;
	assign phi_42__fork_4__valid__0__anchor__out = phi_42_out1_valid;
	assign phi_42_out1_ready = phi_42__fork_4__ready__0__anchor__in;
	assign phi_42__fork_4__ready__0__anchor__out = fork_4_in1_ready;
	assign cst_10_clk = clk;
	assign cst_10_rst = rst;
	assign shl_43_in2_data = cst_10__shl_43__data__0__anchor__in;
	assign cst_10__shl_43__data__0__anchor__out = cst_10_out1_data;
	assign shl_43_in2_valid = cst_10__shl_43__valid__0__anchor__in;
	assign cst_10__shl_43__valid__0__anchor__out = cst_10_out1_valid;
	assign cst_10_out1_ready = cst_10__shl_43__ready__0__anchor__in;
	assign cst_10__shl_43__ready__0__anchor__out = shl_43_in2_ready;
	assign shl_43_clk = clk;
	assign shl_43_rst = rst;
	assign add_44_in1_data = shl_43__add_44__data__0__anchor__in;
	assign shl_43__add_44__data__0__anchor__out = shl_43_out1_data;
	assign add_44_in1_valid = shl_43__add_44__valid__0__anchor__in;
	assign shl_43__add_44__valid__0__anchor__out = shl_43_out1_valid;
	assign shl_43_out1_ready = shl_43__add_44__ready__0__anchor__in;
	assign shl_43__add_44__ready__0__anchor__out = add_44_in1_ready;
	assign add_44_clk = clk;
	assign add_44_rst = rst;
	assign load_47_in2_data = add_44__load_47__data__0__anchor__in;
	assign add_44__load_47__data__0__anchor__out = add_44_out1_data;
	assign load_47_in2_valid = add_44__load_47__valid__0__anchor__in;
	assign add_44__load_47__valid__0__anchor__out = add_44_out1_valid;
	assign add_44_out1_ready = add_44__load_47__ready__0__anchor__in;
	assign add_44__load_47__ready__0__anchor__out = load_47_in2_ready;
	assign load_47_clk = clk;
	assign load_47_rst = rst;
	assign mul_48_in1_data = load_47__mul_48__data__0__anchor__in;
	assign load_47__mul_48__data__0__anchor__out = load_47_out1_data;
	assign mul_48_in1_valid = load_47__mul_48__valid__0__anchor__in;
	assign load_47__mul_48__valid__0__anchor__out = load_47_out1_valid;
	assign load_47_out1_ready = load_47__mul_48__ready__0__anchor__in;
	assign load_47__mul_48__ready__0__anchor__out = mul_48_in1_ready;
	assign MC_A_in5_data = load_47__MC_A__data__0__anchor__in;
	assign load_47__MC_A__data__0__anchor__out = load_47_out2_data;
	assign MC_A_in5_valid = load_47__MC_A__valid__0__anchor__in;
	assign load_47__MC_A__valid__0__anchor__out = load_47_out2_valid;
	assign load_47_out2_ready = load_47__MC_A__ready__0__anchor__in;
	assign load_47__MC_A__ready__0__anchor__out = MC_A_in5_ready;
	assign mul_48_clk = clk;
	assign mul_48_rst = rst;
	assign mul_52_in1_data = mul_48__mul_52__data__0__anchor__in;
	assign mul_48__mul_52__data__0__anchor__out = mul_48_out1_data;
	assign mul_52_in1_valid = mul_48__mul_52__valid__0__anchor__in;
	assign mul_48__mul_52__valid__0__anchor__out = mul_48_out1_valid;
	assign mul_48_out1_ready = mul_48__mul_52__ready__0__anchor__in;
	assign mul_48__mul_52__ready__0__anchor__out = mul_52_in1_ready;
	assign load_51_clk = clk;
	assign load_51_rst = rst;
	assign mul_52_in2_data = load_51__mul_52__data__0__anchor__in;
	assign load_51__mul_52__data__0__anchor__out = load_51_out1_data;
	assign mul_52_in2_valid = load_51__mul_52__valid__0__anchor__in;
	assign load_51__mul_52__valid__0__anchor__out = load_51_out1_valid;
	assign load_51_out1_ready = load_51__mul_52__ready__0__anchor__in;
	assign load_51__mul_52__ready__0__anchor__out = mul_52_in2_ready;
	assign MC_y_in1_data = load_51__MC_y__data__0__anchor__in;
	assign load_51__MC_y__data__0__anchor__out = load_51_out2_data;
	assign MC_y_in1_valid = load_51__MC_y__valid__0__anchor__in;
	assign load_51__MC_y__valid__0__anchor__out = load_51_out2_valid;
	assign load_51_out2_ready = load_51__MC_y__ready__0__anchor__in;
	assign load_51__MC_y__ready__0__anchor__out = MC_y_in1_ready;
	assign mul_52_clk = clk;
	assign mul_52_rst = rst;
	assign add_53_in2_data = mul_52__add_53__data__0__anchor__in;
	assign mul_52__add_53__data__0__anchor__out = mul_52_out1_data;
	assign add_53_in2_valid = mul_52__add_53__valid__0__anchor__in;
	assign mul_52__add_53__valid__0__anchor__out = mul_52_out1_valid;
	assign mul_52_out1_ready = mul_52__add_53__ready__0__anchor__in;
	assign mul_52__add_53__ready__0__anchor__out = add_53_in2_ready;
	assign add_53_clk = clk;
	assign add_53_rst = rst;
	assign branch_22_in1_data = add_53__branch_22__data__0__anchor__in;
	assign add_53__branch_22__data__0__anchor__out = add_53_out1_data;
	assign branch_22_in1_valid = add_53__branch_22__valid__0__anchor__in;
	assign add_53__branch_22__valid__0__anchor__out = add_53_out1_valid;
	assign add_53_out1_ready = add_53__branch_22__ready__0__anchor__in;
	assign add_53__branch_22__ready__0__anchor__out = branch_22_in1_ready;
	assign cst_11_clk = clk;
	assign cst_11_rst = rst;
	assign add_54_in2_data = cst_11__add_54__data__0__anchor__in;
	assign cst_11__add_54__data__0__anchor__out = cst_11_out1_data;
	assign add_54_in2_valid = cst_11__add_54__valid__0__anchor__in;
	assign cst_11__add_54__valid__0__anchor__out = cst_11_out1_valid;
	assign cst_11_out1_ready = cst_11__add_54__ready__0__anchor__in;
	assign cst_11__add_54__ready__0__anchor__out = add_54_in2_ready;
	assign add_54_clk = clk;
	assign add_54_rst = rst;
	assign fork_6_in1_data = add_54__fork_6__data__0__anchor__in;
	assign add_54__fork_6__data__0__anchor__out = add_54_out1_data;
	assign fork_6_in1_valid = add_54__fork_6__valid__0__anchor__in;
	assign add_54__fork_6__valid__0__anchor__out = add_54_out1_valid;
	assign add_54_out1_ready = add_54__fork_6__ready__0__anchor__in;
	assign add_54__fork_6__ready__0__anchor__out = fork_6_in1_ready;
	assign cst_12_clk = clk;
	assign cst_12_rst = rst;
	assign icmp_55_in2_data = cst_12__icmp_55__data__0__anchor__in;
	assign cst_12__icmp_55__data__0__anchor__out = cst_12_out1_data;
	assign icmp_55_in2_valid = cst_12__icmp_55__valid__0__anchor__in;
	assign cst_12__icmp_55__valid__0__anchor__out = cst_12_out1_valid;
	assign cst_12_out1_ready = cst_12__icmp_55__ready__0__anchor__in;
	assign cst_12__icmp_55__ready__0__anchor__out = icmp_55_in2_ready;
	assign icmp_55_clk = clk;
	assign icmp_55_rst = rst;
	assign fork_35_in1_data = icmp_55__fork_35__data__0__anchor__in;
	assign icmp_55__fork_35__data__0__anchor__out = icmp_55_out1_data;
	assign fork_35_in1_valid = icmp_55__fork_35__valid__0__anchor__in;
	assign icmp_55__fork_35__valid__0__anchor__out = icmp_55_out1_valid;
	assign icmp_55_out1_ready = icmp_55__fork_35__ready__0__anchor__in;
	assign icmp_55__fork_35__ready__0__anchor__out = fork_35_in1_ready;
	assign store_1_clk = clk;
	assign store_1_rst = rst;
	assign MC_x_in5_data = store_1__MC_x__data__0__anchor__in;
	assign store_1__MC_x__data__0__anchor__out = store_1_out1_data;
	assign MC_x_in5_valid = store_1__MC_x__valid__0__anchor__in;
	assign store_1__MC_x__valid__0__anchor__out = store_1_out1_valid;
	assign store_1_out1_ready = store_1__MC_x__ready__0__anchor__in;
	assign store_1__MC_x__ready__0__anchor__out = MC_x_in5_ready;
	assign MC_x_in4_data = store_1__MC_x__data__1__anchor__in;
	assign store_1__MC_x__data__1__anchor__out = store_1_out2_data;
	assign MC_x_in4_valid = store_1__MC_x__valid__1__anchor__in;
	assign store_1__MC_x__valid__1__anchor__out = store_1_out2_valid;
	assign store_1_out2_ready = store_1__MC_x__ready__1__anchor__in;
	assign store_1__MC_x__ready__1__anchor__out = MC_x_in4_ready;
	assign cst_13_clk = clk;
	assign cst_13_rst = rst;
	assign add_59_in2_data = cst_13__add_59__data__0__anchor__in;
	assign cst_13__add_59__data__0__anchor__out = cst_13_out1_data;
	assign add_59_in2_valid = cst_13__add_59__valid__0__anchor__in;
	assign cst_13__add_59__valid__0__anchor__out = cst_13_out1_valid;
	assign cst_13_out1_ready = cst_13__add_59__ready__0__anchor__in;
	assign cst_13__add_59__ready__0__anchor__out = add_59_in2_ready;
	assign add_59_clk = clk;
	assign add_59_rst = rst;
	assign fork_7_in1_data = add_59__fork_7__data__0__anchor__in;
	assign add_59__fork_7__data__0__anchor__out = add_59_out1_data;
	assign fork_7_in1_valid = add_59__fork_7__valid__0__anchor__in;
	assign add_59__fork_7__valid__0__anchor__out = add_59_out1_valid;
	assign add_59_out1_ready = add_59__fork_7__ready__0__anchor__in;
	assign add_59__fork_7__ready__0__anchor__out = fork_7_in1_ready;
	assign cst_14_clk = clk;
	assign cst_14_rst = rst;
	assign icmp_60_in2_data = cst_14__icmp_60__data__0__anchor__in;
	assign cst_14__icmp_60__data__0__anchor__out = cst_14_out1_data;
	assign icmp_60_in2_valid = cst_14__icmp_60__valid__0__anchor__in;
	assign cst_14__icmp_60__valid__0__anchor__out = cst_14_out1_valid;
	assign cst_14_out1_ready = cst_14__icmp_60__ready__0__anchor__in;
	assign cst_14__icmp_60__ready__0__anchor__out = icmp_60_in2_ready;
	assign icmp_60_clk = clk;
	assign icmp_60_rst = rst;
	assign fork_36_in1_data = icmp_60__fork_36__data__0__anchor__in;
	assign icmp_60__fork_36__data__0__anchor__out = icmp_60_out1_data;
	assign fork_36_in1_valid = icmp_60__fork_36__valid__0__anchor__in;
	assign icmp_60__fork_36__valid__0__anchor__out = icmp_60_out1_valid;
	assign icmp_60_out1_ready = icmp_60__fork_36__ready__0__anchor__in;
	assign icmp_60__fork_36__ready__0__anchor__out = fork_36_in1_ready;
	assign brCst_block9_clk = clk;
	assign brCst_block9_rst = rst;
	assign fork_37_in1_data = brCst_block9__fork_37__data__0__anchor__in;
	assign brCst_block9__fork_37__data__0__anchor__out = brCst_block9_out1_data;
	assign fork_37_in1_valid = brCst_block9__fork_37__valid__0__anchor__in;
	assign brCst_block9__fork_37__valid__0__anchor__out = brCst_block9_out1_valid;
	assign brCst_block9_out1_ready = brCst_block9__fork_37__ready__0__anchor__in;
	assign brCst_block9__fork_37__ready__0__anchor__out = fork_37_in1_ready;
	assign cst_15_clk = clk;
	assign cst_15_rst = rst;
	assign branch_30_in1_data = cst_15__branch_30__data__0__anchor__in;
	assign cst_15__branch_30__data__0__anchor__out = cst_15_out1_data;
	assign branch_30_in1_valid = cst_15__branch_30__valid__0__anchor__in;
	assign cst_15__branch_30__valid__0__anchor__out = cst_15_out1_valid;
	assign cst_15_out1_ready = cst_15__branch_30__ready__0__anchor__in;
	assign cst_15__branch_30__ready__0__anchor__out = branch_30_in1_ready;
	assign phi_63_clk = clk;
	assign phi_63_rst = rst;
	assign fork_8_in1_data = phi_63__fork_8__data__0__anchor__in;
	assign phi_63__fork_8__data__0__anchor__out = phi_63_out1_data;
	assign fork_8_in1_valid = phi_63__fork_8__valid__0__anchor__in;
	assign phi_63__fork_8__valid__0__anchor__out = phi_63_out1_valid;
	assign phi_63_out1_ready = phi_63__fork_8__ready__0__anchor__in;
	assign phi_63__fork_8__ready__0__anchor__out = fork_8_in1_ready;
	assign load_66_clk = clk;
	assign load_66_rst = rst;
	assign add_70_in1_data = load_66__add_70__data__0__anchor__in;
	assign load_66__add_70__data__0__anchor__out = load_66_out1_data;
	assign add_70_in1_valid = load_66__add_70__valid__0__anchor__in;
	assign load_66__add_70__valid__0__anchor__out = load_66_out1_valid;
	assign load_66_out1_ready = load_66__add_70__ready__0__anchor__in;
	assign load_66__add_70__ready__0__anchor__out = add_70_in1_ready;
	assign MC_x_in6_data = load_66__MC_x__data__0__anchor__in;
	assign load_66__MC_x__data__0__anchor__out = load_66_out2_data;
	assign MC_x_in6_valid = load_66__MC_x__valid__0__anchor__in;
	assign load_66__MC_x__valid__0__anchor__out = load_66_out2_valid;
	assign load_66_out2_ready = load_66__MC_x__ready__0__anchor__in;
	assign load_66__MC_x__ready__0__anchor__out = MC_x_in6_ready;
	assign load_69_clk = clk;
	assign load_69_rst = rst;
	assign add_70_in2_data = load_69__add_70__data__0__anchor__in;
	assign load_69__add_70__data__0__anchor__out = load_69_out1_data;
	assign add_70_in2_valid = load_69__add_70__valid__0__anchor__in;
	assign load_69__add_70__valid__0__anchor__out = load_69_out1_valid;
	assign load_69_out1_ready = load_69__add_70__ready__0__anchor__in;
	assign load_69__add_70__ready__0__anchor__out = add_70_in2_ready;
	assign MC_z_in1_data = load_69__MC_z__data__0__anchor__in;
	assign load_69__MC_z__data__0__anchor__out = load_69_out2_data;
	assign MC_z_in1_valid = load_69__MC_z__valid__0__anchor__in;
	assign load_69__MC_z__valid__0__anchor__out = load_69_out2_valid;
	assign load_69_out2_ready = load_69__MC_z__ready__0__anchor__in;
	assign load_69__MC_z__ready__0__anchor__out = MC_z_in1_ready;
	assign add_70_clk = clk;
	assign add_70_rst = rst;
	assign store_2_in1_data = add_70__store_2__data__0__anchor__in;
	assign add_70__store_2__data__0__anchor__out = add_70_out1_data;
	assign store_2_in1_valid = add_70__store_2__valid__0__anchor__in;
	assign add_70__store_2__valid__0__anchor__out = add_70_out1_valid;
	assign add_70_out1_ready = add_70__store_2__ready__0__anchor__in;
	assign add_70__store_2__ready__0__anchor__out = store_2_in1_ready;
	assign store_2_clk = clk;
	assign store_2_rst = rst;
	assign MC_x_in8_data = store_2__MC_x__data__0__anchor__in;
	assign store_2__MC_x__data__0__anchor__out = store_2_out1_data;
	assign MC_x_in8_valid = store_2__MC_x__valid__0__anchor__in;
	assign store_2__MC_x__valid__0__anchor__out = store_2_out1_valid;
	assign store_2_out1_ready = store_2__MC_x__ready__0__anchor__in;
	assign store_2__MC_x__ready__0__anchor__out = MC_x_in8_ready;
	assign MC_x_in7_data = store_2__MC_x__data__1__anchor__in;
	assign store_2__MC_x__data__1__anchor__out = store_2_out2_data;
	assign MC_x_in7_valid = store_2__MC_x__valid__1__anchor__in;
	assign store_2__MC_x__valid__1__anchor__out = store_2_out2_valid;
	assign store_2_out2_ready = store_2__MC_x__ready__1__anchor__in;
	assign store_2__MC_x__ready__1__anchor__out = MC_x_in7_ready;
	assign cst_16_clk = clk;
	assign cst_16_rst = rst;
	assign add_73_in2_data = cst_16__add_73__data__0__anchor__in;
	assign cst_16__add_73__data__0__anchor__out = cst_16_out1_data;
	assign add_73_in2_valid = cst_16__add_73__valid__0__anchor__in;
	assign cst_16__add_73__valid__0__anchor__out = cst_16_out1_valid;
	assign cst_16_out1_ready = cst_16__add_73__ready__0__anchor__in;
	assign cst_16__add_73__ready__0__anchor__out = add_73_in2_ready;
	assign add_73_clk = clk;
	assign add_73_rst = rst;
	assign fork_9_in1_data = add_73__fork_9__data__0__anchor__in;
	assign add_73__fork_9__data__0__anchor__out = add_73_out1_data;
	assign fork_9_in1_valid = add_73__fork_9__valid__0__anchor__in;
	assign add_73__fork_9__valid__0__anchor__out = add_73_out1_valid;
	assign add_73_out1_ready = add_73__fork_9__ready__0__anchor__in;
	assign add_73__fork_9__ready__0__anchor__out = fork_9_in1_ready;
	assign cst_17_clk = clk;
	assign cst_17_rst = rst;
	assign icmp_74_in2_data = cst_17__icmp_74__data__0__anchor__in;
	assign cst_17__icmp_74__data__0__anchor__out = cst_17_out1_data;
	assign icmp_74_in2_valid = cst_17__icmp_74__valid__0__anchor__in;
	assign cst_17__icmp_74__valid__0__anchor__out = cst_17_out1_valid;
	assign cst_17_out1_ready = cst_17__icmp_74__ready__0__anchor__in;
	assign cst_17__icmp_74__ready__0__anchor__out = icmp_74_in2_ready;
	assign icmp_74_clk = clk;
	assign icmp_74_rst = rst;
	assign fork_38_in1_data = icmp_74__fork_38__data__0__anchor__in;
	assign icmp_74__fork_38__data__0__anchor__out = icmp_74_out1_data;
	assign fork_38_in1_valid = icmp_74__fork_38__valid__0__anchor__in;
	assign icmp_74__fork_38__valid__0__anchor__out = icmp_74_out1_valid;
	assign icmp_74_out1_ready = icmp_74__fork_38__ready__0__anchor__in;
	assign icmp_74__fork_38__ready__0__anchor__out = fork_38_in1_ready;
	assign brCst_block11_clk = clk;
	assign brCst_block11_rst = rst;
	assign fork_39_in1_data = brCst_block11__fork_39__data__0__anchor__in;
	assign brCst_block11__fork_39__data__0__anchor__out = brCst_block11_out1_data;
	assign fork_39_in1_valid = brCst_block11__fork_39__valid__0__anchor__in;
	assign brCst_block11__fork_39__valid__0__anchor__out = brCst_block11_out1_valid;
	assign brCst_block11_out1_ready = brCst_block11__fork_39__ready__0__anchor__in;
	assign brCst_block11__fork_39__ready__0__anchor__out = fork_39_in1_ready;
	assign cst_18_clk = clk;
	assign cst_18_rst = rst;
	assign branch_34_in1_data = cst_18__branch_34__data__0__anchor__in;
	assign cst_18__branch_34__data__0__anchor__out = cst_18_out1_data;
	assign branch_34_in1_valid = cst_18__branch_34__valid__0__anchor__in;
	assign cst_18__branch_34__valid__0__anchor__out = cst_18_out1_valid;
	assign cst_18_out1_ready = cst_18__branch_34__ready__0__anchor__in;
	assign cst_18__branch_34__ready__0__anchor__out = branch_34_in1_ready;
	assign phi_77_clk = clk;
	assign phi_77_rst = rst;
	assign fork_10_in1_data = phi_77__fork_10__data__0__anchor__in;
	assign phi_77__fork_10__data__0__anchor__out = phi_77_out1_data;
	assign fork_10_in1_valid = phi_77__fork_10__valid__0__anchor__in;
	assign phi_77__fork_10__valid__0__anchor__out = phi_77_out1_valid;
	assign phi_77_out1_ready = phi_77__fork_10__ready__0__anchor__in;
	assign phi_77__fork_10__ready__0__anchor__out = fork_10_in1_ready;
	assign load_80_clk = clk;
	assign load_80_rst = rst;
	assign branch_36_in1_data = load_80__branch_36__data__0__anchor__in;
	assign load_80__branch_36__data__0__anchor__out = load_80_out1_data;
	assign branch_36_in1_valid = load_80__branch_36__valid__0__anchor__in;
	assign load_80__branch_36__valid__0__anchor__out = load_80_out1_valid;
	assign load_80_out1_ready = load_80__branch_36__ready__0__anchor__in;
	assign load_80__branch_36__ready__0__anchor__out = branch_36_in1_ready;
	assign MC_w_in2_data = load_80__MC_w__data__0__anchor__in;
	assign load_80__MC_w__data__0__anchor__out = load_80_out2_data;
	assign MC_w_in2_valid = load_80__MC_w__valid__0__anchor__in;
	assign load_80__MC_w__valid__0__anchor__out = load_80_out2_valid;
	assign load_80_out2_ready = load_80__MC_w__ready__0__anchor__in;
	assign load_80__MC_w__ready__0__anchor__out = MC_w_in2_ready;
	assign brCst_block12_clk = clk;
	assign brCst_block12_rst = rst;
	assign fork_40_in1_data = brCst_block12__fork_40__data__0__anchor__in;
	assign brCst_block12__fork_40__data__0__anchor__out = brCst_block12_out1_data;
	assign fork_40_in1_valid = brCst_block12__fork_40__valid__0__anchor__in;
	assign brCst_block12__fork_40__valid__0__anchor__out = brCst_block12_out1_valid;
	assign brCst_block12_out1_ready = brCst_block12__fork_40__ready__0__anchor__in;
	assign brCst_block12__fork_40__ready__0__anchor__out = fork_40_in1_ready;
	assign phi_82_clk = clk;
	assign phi_82_rst = rst;
	assign add_94_in1_data = phi_82__add_94__data__0__anchor__in;
	assign phi_82__add_94__data__0__anchor__out = phi_82_out1_data;
	assign add_94_in1_valid = phi_82__add_94__valid__0__anchor__in;
	assign phi_82__add_94__valid__0__anchor__out = phi_82_out1_valid;
	assign phi_82_out1_ready = phi_82__add_94__ready__0__anchor__in;
	assign phi_82__add_94__ready__0__anchor__out = add_94_in1_ready;
	assign cst_19_clk = clk;
	assign cst_19_rst = rst;
	assign branch_37_in1_data = cst_19__branch_37__data__0__anchor__in;
	assign cst_19__branch_37__data__0__anchor__out = cst_19_out1_data;
	assign branch_37_in1_valid = cst_19__branch_37__valid__0__anchor__in;
	assign cst_19__branch_37__valid__0__anchor__out = cst_19_out1_valid;
	assign cst_19_out1_ready = cst_19__branch_37__ready__0__anchor__in;
	assign cst_19__branch_37__ready__0__anchor__out = branch_37_in1_ready;
	assign phi_83_clk = clk;
	assign phi_83_rst = rst;
	assign fork_11_in1_data = phi_83__fork_11__data__0__anchor__in;
	assign phi_83__fork_11__data__0__anchor__out = phi_83_out1_data;
	assign fork_11_in1_valid = phi_83__fork_11__valid__0__anchor__in;
	assign phi_83__fork_11__valid__0__anchor__out = phi_83_out1_valid;
	assign phi_83_out1_ready = phi_83__fork_11__ready__0__anchor__in;
	assign phi_83__fork_11__ready__0__anchor__out = fork_11_in1_ready;
	assign cst_20_clk = clk;
	assign cst_20_rst = rst;
	assign shl_84_in2_data = cst_20__shl_84__data__0__anchor__in;
	assign cst_20__shl_84__data__0__anchor__out = cst_20_out1_data;
	assign shl_84_in2_valid = cst_20__shl_84__valid__0__anchor__in;
	assign cst_20__shl_84__valid__0__anchor__out = cst_20_out1_valid;
	assign cst_20_out1_ready = cst_20__shl_84__ready__0__anchor__in;
	assign cst_20__shl_84__ready__0__anchor__out = shl_84_in2_ready;
	assign shl_84_clk = clk;
	assign shl_84_rst = rst;
	assign add_85_in1_data = shl_84__add_85__data__0__anchor__in;
	assign shl_84__add_85__data__0__anchor__out = shl_84_out1_data;
	assign add_85_in1_valid = shl_84__add_85__valid__0__anchor__in;
	assign shl_84__add_85__valid__0__anchor__out = shl_84_out1_valid;
	assign shl_84_out1_ready = shl_84__add_85__ready__0__anchor__in;
	assign shl_84__add_85__ready__0__anchor__out = add_85_in1_ready;
	assign add_85_clk = clk;
	assign add_85_rst = rst;
	assign load_88_in2_data = add_85__load_88__data__0__anchor__in;
	assign add_85__load_88__data__0__anchor__out = add_85_out1_data;
	assign load_88_in2_valid = add_85__load_88__valid__0__anchor__in;
	assign add_85__load_88__valid__0__anchor__out = add_85_out1_valid;
	assign add_85_out1_ready = add_85__load_88__ready__0__anchor__in;
	assign add_85__load_88__ready__0__anchor__out = load_88_in2_ready;
	assign load_88_clk = clk;
	assign load_88_rst = rst;
	assign mul_89_in1_data = load_88__mul_89__data__0__anchor__in;
	assign load_88__mul_89__data__0__anchor__out = load_88_out1_data;
	assign mul_89_in1_valid = load_88__mul_89__valid__0__anchor__in;
	assign load_88__mul_89__valid__0__anchor__out = load_88_out1_valid;
	assign load_88_out1_ready = load_88__mul_89__ready__0__anchor__in;
	assign load_88__mul_89__ready__0__anchor__out = mul_89_in1_ready;
	assign MC_A_in6_data = load_88__MC_A__data__0__anchor__in;
	assign load_88__MC_A__data__0__anchor__out = load_88_out2_data;
	assign MC_A_in6_valid = load_88__MC_A__valid__0__anchor__in;
	assign load_88__MC_A__valid__0__anchor__out = load_88_out2_valid;
	assign load_88_out2_ready = load_88__MC_A__ready__0__anchor__in;
	assign load_88__MC_A__ready__0__anchor__out = MC_A_in6_ready;
	assign mul_89_clk = clk;
	assign mul_89_rst = rst;
	assign mul_93_in1_data = mul_89__mul_93__data__0__anchor__in;
	assign mul_89__mul_93__data__0__anchor__out = mul_89_out1_data;
	assign mul_93_in1_valid = mul_89__mul_93__valid__0__anchor__in;
	assign mul_89__mul_93__valid__0__anchor__out = mul_89_out1_valid;
	assign mul_89_out1_ready = mul_89__mul_93__ready__0__anchor__in;
	assign mul_89__mul_93__ready__0__anchor__out = mul_93_in1_ready;
	assign load_92_clk = clk;
	assign load_92_rst = rst;
	assign mul_93_in2_data = load_92__mul_93__data__0__anchor__in;
	assign load_92__mul_93__data__0__anchor__out = load_92_out1_data;
	assign mul_93_in2_valid = load_92__mul_93__valid__0__anchor__in;
	assign load_92__mul_93__valid__0__anchor__out = load_92_out1_valid;
	assign load_92_out1_ready = load_92__mul_93__ready__0__anchor__in;
	assign load_92__mul_93__ready__0__anchor__out = mul_93_in2_ready;
	assign MC_x_in9_data = load_92__MC_x__data__0__anchor__in;
	assign load_92__MC_x__data__0__anchor__out = load_92_out2_data;
	assign MC_x_in9_valid = load_92__MC_x__valid__0__anchor__in;
	assign load_92__MC_x__valid__0__anchor__out = load_92_out2_valid;
	assign load_92_out2_ready = load_92__MC_x__ready__0__anchor__in;
	assign load_92__MC_x__ready__0__anchor__out = MC_x_in9_ready;
	assign mul_93_clk = clk;
	assign mul_93_rst = rst;
	assign add_94_in2_data = mul_93__add_94__data__0__anchor__in;
	assign mul_93__add_94__data__0__anchor__out = mul_93_out1_data;
	assign add_94_in2_valid = mul_93__add_94__valid__0__anchor__in;
	assign mul_93__add_94__valid__0__anchor__out = mul_93_out1_valid;
	assign mul_93_out1_ready = mul_93__add_94__ready__0__anchor__in;
	assign mul_93__add_94__ready__0__anchor__out = add_94_in2_ready;
	assign add_94_clk = clk;
	assign add_94_rst = rst;
	assign branch_40_in1_data = add_94__branch_40__data__0__anchor__in;
	assign add_94__branch_40__data__0__anchor__out = add_94_out1_data;
	assign branch_40_in1_valid = add_94__branch_40__valid__0__anchor__in;
	assign add_94__branch_40__valid__0__anchor__out = add_94_out1_valid;
	assign add_94_out1_ready = add_94__branch_40__ready__0__anchor__in;
	assign add_94__branch_40__ready__0__anchor__out = branch_40_in1_ready;
	assign cst_21_clk = clk;
	assign cst_21_rst = rst;
	assign add_95_in2_data = cst_21__add_95__data__0__anchor__in;
	assign cst_21__add_95__data__0__anchor__out = cst_21_out1_data;
	assign add_95_in2_valid = cst_21__add_95__valid__0__anchor__in;
	assign cst_21__add_95__valid__0__anchor__out = cst_21_out1_valid;
	assign cst_21_out1_ready = cst_21__add_95__ready__0__anchor__in;
	assign cst_21__add_95__ready__0__anchor__out = add_95_in2_ready;
	assign add_95_clk = clk;
	assign add_95_rst = rst;
	assign fork_13_in1_data = add_95__fork_13__data__0__anchor__in;
	assign add_95__fork_13__data__0__anchor__out = add_95_out1_data;
	assign fork_13_in1_valid = add_95__fork_13__valid__0__anchor__in;
	assign add_95__fork_13__valid__0__anchor__out = add_95_out1_valid;
	assign add_95_out1_ready = add_95__fork_13__ready__0__anchor__in;
	assign add_95__fork_13__ready__0__anchor__out = fork_13_in1_ready;
	assign cst_22_clk = clk;
	assign cst_22_rst = rst;
	assign icmp_96_in2_data = cst_22__icmp_96__data__0__anchor__in;
	assign cst_22__icmp_96__data__0__anchor__out = cst_22_out1_data;
	assign icmp_96_in2_valid = cst_22__icmp_96__valid__0__anchor__in;
	assign cst_22__icmp_96__valid__0__anchor__out = cst_22_out1_valid;
	assign cst_22_out1_ready = cst_22__icmp_96__ready__0__anchor__in;
	assign cst_22__icmp_96__ready__0__anchor__out = icmp_96_in2_ready;
	assign icmp_96_clk = clk;
	assign icmp_96_rst = rst;
	assign fork_41_in1_data = icmp_96__fork_41__data__0__anchor__in;
	assign icmp_96__fork_41__data__0__anchor__out = icmp_96_out1_data;
	assign fork_41_in1_valid = icmp_96__fork_41__valid__0__anchor__in;
	assign icmp_96__fork_41__valid__0__anchor__out = icmp_96_out1_valid;
	assign icmp_96_out1_ready = icmp_96__fork_41__ready__0__anchor__in;
	assign icmp_96__fork_41__ready__0__anchor__out = fork_41_in1_ready;
	assign store_3_clk = clk;
	assign store_3_rst = rst;
	assign MC_w_in4_data = store_3__MC_w__data__0__anchor__in;
	assign store_3__MC_w__data__0__anchor__out = store_3_out1_data;
	assign MC_w_in4_valid = store_3__MC_w__valid__0__anchor__in;
	assign store_3__MC_w__valid__0__anchor__out = store_3_out1_valid;
	assign store_3_out1_ready = store_3__MC_w__ready__0__anchor__in;
	assign store_3__MC_w__ready__0__anchor__out = MC_w_in4_ready;
	assign MC_w_in3_data = store_3__MC_w__data__1__anchor__in;
	assign store_3__MC_w__data__1__anchor__out = store_3_out2_data;
	assign MC_w_in3_valid = store_3__MC_w__valid__1__anchor__in;
	assign store_3__MC_w__valid__1__anchor__out = store_3_out2_valid;
	assign store_3_out2_ready = store_3__MC_w__ready__1__anchor__in;
	assign store_3__MC_w__ready__1__anchor__out = MC_w_in3_ready;
	assign cst_23_clk = clk;
	assign cst_23_rst = rst;
	assign add_100_in2_data = cst_23__add_100__data__0__anchor__in;
	assign cst_23__add_100__data__0__anchor__out = cst_23_out1_data;
	assign add_100_in2_valid = cst_23__add_100__valid__0__anchor__in;
	assign cst_23__add_100__valid__0__anchor__out = cst_23_out1_valid;
	assign cst_23_out1_ready = cst_23__add_100__ready__0__anchor__in;
	assign cst_23__add_100__ready__0__anchor__out = add_100_in2_ready;
	assign add_100_clk = clk;
	assign add_100_rst = rst;
	assign fork_14_in1_data = add_100__fork_14__data__0__anchor__in;
	assign add_100__fork_14__data__0__anchor__out = add_100_out1_data;
	assign fork_14_in1_valid = add_100__fork_14__valid__0__anchor__in;
	assign add_100__fork_14__valid__0__anchor__out = add_100_out1_valid;
	assign add_100_out1_ready = add_100__fork_14__ready__0__anchor__in;
	assign add_100__fork_14__ready__0__anchor__out = fork_14_in1_ready;
	assign cst_24_clk = clk;
	assign cst_24_rst = rst;
	assign icmp_101_in2_data = cst_24__icmp_101__data__0__anchor__in;
	assign cst_24__icmp_101__data__0__anchor__out = cst_24_out1_data;
	assign icmp_101_in2_valid = cst_24__icmp_101__valid__0__anchor__in;
	assign cst_24__icmp_101__valid__0__anchor__out = cst_24_out1_valid;
	assign cst_24_out1_ready = cst_24__icmp_101__ready__0__anchor__in;
	assign cst_24__icmp_101__ready__0__anchor__out = icmp_101_in2_ready;
	assign icmp_101_clk = clk;
	assign icmp_101_rst = rst;
	assign fork_42_in1_data = icmp_101__fork_42__data__0__anchor__in;
	assign icmp_101__fork_42__data__0__anchor__out = icmp_101_out1_data;
	assign fork_42_in1_valid = icmp_101__fork_42__valid__0__anchor__in;
	assign icmp_101__fork_42__valid__0__anchor__out = icmp_101_out1_valid;
	assign icmp_101_out1_ready = icmp_101__fork_42__ready__0__anchor__in;
	assign icmp_101__fork_42__ready__0__anchor__out = fork_42_in1_ready;
	assign ret_0_clk = clk;
	assign ret_0_rst = rst;
	assign end_0_in10_data = ret_0__end_0__data__0__anchor__in;
	assign ret_0__end_0__data__0__anchor__out = ret_0_out1_data;
	assign end_0_in10_valid = ret_0__end_0__valid__0__anchor__in;
	assign ret_0__end_0__valid__0__anchor__out = ret_0_out1_valid;
	assign ret_0_out1_ready = ret_0__end_0__ready__0__anchor__in;
	assign ret_0__end_0__ready__0__anchor__out = end_0_in10_ready;
	assign phi_n0_clk = clk;
	assign phi_n0_rst = rst;
	assign branch_5_in1_data = phi_n0__branch_5__data__0__anchor__in;
	assign phi_n0__branch_5__data__0__anchor__out = phi_n0_out1_data;
	assign branch_5_in1_valid = phi_n0__branch_5__valid__0__anchor__in;
	assign phi_n0__branch_5__valid__0__anchor__out = phi_n0_out1_valid;
	assign phi_n0_out1_ready = phi_n0__branch_5__ready__0__anchor__in;
	assign phi_n0__branch_5__ready__0__anchor__out = branch_5_in1_ready;
	assign phi_n1_clk = clk;
	assign phi_n1_rst = rst;
	assign branch_6_in1_data = phi_n1__branch_6__data__0__anchor__in;
	assign phi_n1__branch_6__data__0__anchor__out = phi_n1_out1_data;
	assign branch_6_in1_valid = phi_n1__branch_6__valid__0__anchor__in;
	assign phi_n1__branch_6__valid__0__anchor__out = phi_n1_out1_valid;
	assign phi_n1_out1_ready = phi_n1__branch_6__ready__0__anchor__in;
	assign phi_n1__branch_6__ready__0__anchor__out = branch_6_in1_ready;
	assign phi_n2_clk = clk;
	assign phi_n2_rst = rst;
	assign add_32_in1_data = phi_n2__add_32__data__0__anchor__in;
	assign phi_n2__add_32__data__0__anchor__out = phi_n2_out1_data;
	assign add_32_in1_valid = phi_n2__add_32__valid__0__anchor__in;
	assign phi_n2__add_32__valid__0__anchor__out = phi_n2_out1_valid;
	assign phi_n2_out1_ready = phi_n2__add_32__ready__0__anchor__in;
	assign phi_n2__add_32__ready__0__anchor__out = add_32_in1_ready;
	assign phi_n3_clk = clk;
	assign phi_n3_rst = rst;
	assign branch_12_in1_data = phi_n3__branch_12__data__0__anchor__in;
	assign phi_n3__branch_12__data__0__anchor__out = phi_n3_out1_data;
	assign branch_12_in1_valid = phi_n3__branch_12__valid__0__anchor__in;
	assign phi_n3__branch_12__valid__0__anchor__out = phi_n3_out1_valid;
	assign phi_n3_out1_ready = phi_n3__branch_12__ready__0__anchor__in;
	assign phi_n3__branch_12__ready__0__anchor__out = branch_12_in1_ready;
	assign phi_n4_clk = clk;
	assign phi_n4_rst = rst;
	assign branch_13_in1_data = phi_n4__branch_13__data__0__anchor__in;
	assign phi_n4__branch_13__data__0__anchor__out = phi_n4_out1_data;
	assign branch_13_in1_valid = phi_n4__branch_13__valid__0__anchor__in;
	assign phi_n4__branch_13__valid__0__anchor__out = phi_n4_out1_valid;
	assign phi_n4_out1_ready = phi_n4__branch_13__ready__0__anchor__in;
	assign phi_n4__branch_13__ready__0__anchor__out = branch_13_in1_ready;
	assign phi_n5_clk = clk;
	assign phi_n5_rst = rst;
	assign fork_17_in1_data = phi_n5__fork_17__data__0__anchor__in;
	assign phi_n5__fork_17__data__0__anchor__out = phi_n5_out1_data;
	assign fork_17_in1_valid = phi_n5__fork_17__valid__0__anchor__in;
	assign phi_n5__fork_17__valid__0__anchor__out = phi_n5_out1_valid;
	assign phi_n5_out1_ready = phi_n5__fork_17__ready__0__anchor__in;
	assign phi_n5__fork_17__ready__0__anchor__out = fork_17_in1_ready;
	assign phi_n6_clk = clk;
	assign phi_n6_rst = rst;
	assign branch_9_in1_data = phi_n6__branch_9__data__0__anchor__in;
	assign phi_n6__branch_9__data__0__anchor__out = phi_n6_out1_data;
	assign branch_9_in1_valid = phi_n6__branch_9__valid__0__anchor__in;
	assign phi_n6__branch_9__valid__0__anchor__out = phi_n6_out1_valid;
	assign phi_n6_out1_ready = phi_n6__branch_9__ready__0__anchor__in;
	assign phi_n6__branch_9__ready__0__anchor__out = branch_9_in1_ready;
	assign phi_n7_clk = clk;
	assign phi_n7_rst = rst;
	assign branch_10_in1_data = phi_n7__branch_10__data__0__anchor__in;
	assign phi_n7__branch_10__data__0__anchor__out = phi_n7_out1_data;
	assign branch_10_in1_valid = phi_n7__branch_10__valid__0__anchor__in;
	assign phi_n7__branch_10__valid__0__anchor__out = phi_n7_out1_valid;
	assign phi_n7_out1_ready = phi_n7__branch_10__ready__0__anchor__in;
	assign phi_n7__branch_10__ready__0__anchor__out = branch_10_in1_ready;
	assign phi_n8_clk = clk;
	assign phi_n8_rst = rst;
	assign branch_15_in1_data = phi_n8__branch_15__data__0__anchor__in;
	assign phi_n8__branch_15__data__0__anchor__out = phi_n8_out1_data;
	assign branch_15_in1_valid = phi_n8__branch_15__valid__0__anchor__in;
	assign phi_n8__branch_15__valid__0__anchor__out = phi_n8_out1_valid;
	assign phi_n8_out1_ready = phi_n8__branch_15__ready__0__anchor__in;
	assign phi_n8__branch_15__ready__0__anchor__out = branch_15_in1_ready;
	assign phi_n9_clk = clk;
	assign phi_n9_rst = rst;
	assign branch_16_in1_data = phi_n9__branch_16__data__0__anchor__in;
	assign phi_n9__branch_16__data__0__anchor__out = phi_n9_out1_data;
	assign branch_16_in1_valid = phi_n9__branch_16__valid__0__anchor__in;
	assign phi_n9__branch_16__valid__0__anchor__out = phi_n9_out1_valid;
	assign phi_n9_out1_ready = phi_n9__branch_16__ready__0__anchor__in;
	assign phi_n9__branch_16__ready__0__anchor__out = branch_16_in1_ready;
	assign phi_n10_clk = clk;
	assign phi_n10_rst = rst;
	assign branch_19_in1_data = phi_n10__branch_19__data__0__anchor__in;
	assign phi_n10__branch_19__data__0__anchor__out = phi_n10_out1_data;
	assign branch_19_in1_valid = phi_n10__branch_19__valid__0__anchor__in;
	assign phi_n10__branch_19__valid__0__anchor__out = phi_n10_out1_valid;
	assign phi_n10_out1_ready = phi_n10__branch_19__ready__0__anchor__in;
	assign phi_n10__branch_19__ready__0__anchor__out = branch_19_in1_ready;
	assign phi_n11_clk = clk;
	assign phi_n11_rst = rst;
	assign branch_20_in1_data = phi_n11__branch_20__data__0__anchor__in;
	assign phi_n11__branch_20__data__0__anchor__out = phi_n11_out1_data;
	assign branch_20_in1_valid = phi_n11__branch_20__valid__0__anchor__in;
	assign phi_n11__branch_20__valid__0__anchor__out = phi_n11_out1_valid;
	assign phi_n11_out1_ready = phi_n11__branch_20__ready__0__anchor__in;
	assign phi_n11__branch_20__ready__0__anchor__out = branch_20_in1_ready;
	assign phi_n12_clk = clk;
	assign phi_n12_rst = rst;
	assign store_1_in1_data = phi_n12__store_1__data__0__anchor__in;
	assign phi_n12__store_1__data__0__anchor__out = phi_n12_out1_data;
	assign store_1_in1_valid = phi_n12__store_1__valid__0__anchor__in;
	assign phi_n12__store_1__valid__0__anchor__out = phi_n12_out1_valid;
	assign phi_n12_out1_ready = phi_n12__store_1__ready__0__anchor__in;
	assign phi_n12__store_1__ready__0__anchor__out = store_1_in1_ready;
	assign phi_n13_clk = clk;
	assign phi_n13_rst = rst;
	assign fork_20_in1_data = phi_n13__fork_20__data__0__anchor__in;
	assign phi_n13__fork_20__data__0__anchor__out = phi_n13_out1_data;
	assign fork_20_in1_valid = phi_n13__fork_20__valid__0__anchor__in;
	assign phi_n13__fork_20__valid__0__anchor__out = phi_n13_out1_valid;
	assign phi_n13_out1_ready = phi_n13__fork_20__ready__0__anchor__in;
	assign phi_n13__fork_20__ready__0__anchor__out = fork_20_in1_ready;
	assign phi_n14_clk = clk;
	assign phi_n14_rst = rst;
	assign branch_27_in1_data = phi_n14__branch_27__data__0__anchor__in;
	assign phi_n14__branch_27__data__0__anchor__out = phi_n14_out1_data;
	assign branch_27_in1_valid = phi_n14__branch_27__valid__0__anchor__in;
	assign phi_n14__branch_27__valid__0__anchor__out = phi_n14_out1_valid;
	assign phi_n14_out1_ready = phi_n14__branch_27__ready__0__anchor__in;
	assign phi_n14__branch_27__ready__0__anchor__out = branch_27_in1_ready;
	assign phi_n15_clk = clk;
	assign phi_n15_rst = rst;
	assign branch_29_in1_data = phi_n15__branch_29__data__0__anchor__in;
	assign phi_n15__branch_29__data__0__anchor__out = phi_n15_out1_data;
	assign branch_29_in1_valid = phi_n15__branch_29__valid__0__anchor__in;
	assign phi_n15__branch_29__valid__0__anchor__out = phi_n15_out1_valid;
	assign phi_n15_out1_ready = phi_n15__branch_29__ready__0__anchor__in;
	assign phi_n15__branch_29__ready__0__anchor__out = branch_29_in1_ready;
	assign phi_n16_clk = clk;
	assign phi_n16_rst = rst;
	assign fork_22_in1_data = phi_n16__fork_22__data__0__anchor__in;
	assign phi_n16__fork_22__data__0__anchor__out = phi_n16_out1_data;
	assign fork_22_in1_valid = phi_n16__fork_22__valid__0__anchor__in;
	assign phi_n16__fork_22__valid__0__anchor__out = phi_n16_out1_valid;
	assign phi_n16_out1_ready = phi_n16__fork_22__ready__0__anchor__in;
	assign phi_n16__fork_22__ready__0__anchor__out = fork_22_in1_ready;
	assign phi_n17_clk = clk;
	assign phi_n17_rst = rst;
	assign fork_23_in1_data = phi_n17__fork_23__data__0__anchor__in;
	assign phi_n17__fork_23__data__0__anchor__out = phi_n17_out1_data;
	assign fork_23_in1_valid = phi_n17__fork_23__valid__0__anchor__in;
	assign phi_n17__fork_23__valid__0__anchor__out = phi_n17_out1_valid;
	assign phi_n17_out1_ready = phi_n17__fork_23__ready__0__anchor__in;
	assign phi_n17__fork_23__ready__0__anchor__out = fork_23_in1_ready;
	assign phi_n18_clk = clk;
	assign phi_n18_rst = rst;
	assign branch_26_in1_data = phi_n18__branch_26__data__0__anchor__in;
	assign phi_n18__branch_26__data__0__anchor__out = phi_n18_out1_data;
	assign branch_26_in1_valid = phi_n18__branch_26__valid__0__anchor__in;
	assign phi_n18__branch_26__valid__0__anchor__out = phi_n18_out1_valid;
	assign phi_n18_out1_ready = phi_n18__branch_26__ready__0__anchor__in;
	assign phi_n18__branch_26__ready__0__anchor__out = branch_26_in1_ready;
	assign phi_n19_clk = clk;
	assign phi_n19_rst = rst;
	assign branch_31_in1_data = phi_n19__branch_31__data__0__anchor__in;
	assign phi_n19__branch_31__data__0__anchor__out = phi_n19_out1_data;
	assign branch_31_in1_valid = phi_n19__branch_31__valid__0__anchor__in;
	assign phi_n19__branch_31__valid__0__anchor__out = phi_n19_out1_valid;
	assign phi_n19_out1_ready = phi_n19__branch_31__ready__0__anchor__in;
	assign phi_n19__branch_31__ready__0__anchor__out = branch_31_in1_ready;
	assign phi_n20_clk = clk;
	assign phi_n20_rst = rst;
	assign branch_33_in1_data = phi_n20__branch_33__data__0__anchor__in;
	assign phi_n20__branch_33__data__0__anchor__out = phi_n20_out1_data;
	assign branch_33_in1_valid = phi_n20__branch_33__valid__0__anchor__in;
	assign phi_n20__branch_33__valid__0__anchor__out = phi_n20_out1_valid;
	assign phi_n20_out1_ready = phi_n20__branch_33__ready__0__anchor__in;
	assign phi_n20__branch_33__ready__0__anchor__out = branch_33_in1_ready;
	assign phi_n21_clk = clk;
	assign phi_n21_rst = rst;
	assign branch_35_in1_data = phi_n21__branch_35__data__0__anchor__in;
	assign phi_n21__branch_35__data__0__anchor__out = phi_n21_out1_data;
	assign branch_35_in1_valid = phi_n21__branch_35__valid__0__anchor__in;
	assign phi_n21__branch_35__valid__0__anchor__out = phi_n21_out1_valid;
	assign phi_n21_out1_ready = phi_n21__branch_35__ready__0__anchor__in;
	assign phi_n21__branch_35__ready__0__anchor__out = branch_35_in1_ready;
	assign phi_n22_clk = clk;
	assign phi_n22_rst = rst;
	assign branch_38_in1_data = phi_n22__branch_38__data__0__anchor__in;
	assign phi_n22__branch_38__data__0__anchor__out = phi_n22_out1_data;
	assign branch_38_in1_valid = phi_n22__branch_38__valid__0__anchor__in;
	assign phi_n22__branch_38__valid__0__anchor__out = phi_n22_out1_valid;
	assign phi_n22_out1_ready = phi_n22__branch_38__ready__0__anchor__in;
	assign phi_n22__branch_38__ready__0__anchor__out = branch_38_in1_ready;
	assign phi_n23_clk = clk;
	assign phi_n23_rst = rst;
	assign store_3_in1_data = phi_n23__store_3__data__0__anchor__in;
	assign phi_n23__store_3__data__0__anchor__out = phi_n23_out1_data;
	assign store_3_in1_valid = phi_n23__store_3__valid__0__anchor__in;
	assign phi_n23__store_3__valid__0__anchor__out = phi_n23_out1_valid;
	assign phi_n23_out1_ready = phi_n23__store_3__ready__0__anchor__in;
	assign phi_n23__store_3__ready__0__anchor__out = store_3_in1_ready;
	assign phi_n24_clk = clk;
	assign phi_n24_rst = rst;
	assign fork_26_in1_data = phi_n24__fork_26__data__0__anchor__in;
	assign phi_n24__fork_26__data__0__anchor__out = phi_n24_out1_data;
	assign fork_26_in1_valid = phi_n24__fork_26__valid__0__anchor__in;
	assign phi_n24__fork_26__valid__0__anchor__out = phi_n24_out1_valid;
	assign phi_n24_out1_ready = phi_n24__fork_26__ready__0__anchor__in;
	assign phi_n24__fork_26__ready__0__anchor__out = fork_26_in1_ready;
	assign phi_n25_clk = clk;
	assign phi_n25_rst = rst;
	assign branch_44_in1_data = phi_n25__branch_44__data__0__anchor__in;
	assign phi_n25__branch_44__data__0__anchor__out = phi_n25_out1_data;
	assign branch_44_in1_valid = phi_n25__branch_44__valid__0__anchor__in;
	assign phi_n25__branch_44__valid__0__anchor__out = phi_n25_out1_valid;
	assign phi_n25_out1_ready = phi_n25__branch_44__ready__0__anchor__in;
	assign phi_n25__branch_44__ready__0__anchor__out = branch_44_in1_ready;
	assign phi_n26_clk = clk;
	assign phi_n26_rst = rst;
	assign fork_27_in1_data = phi_n26__fork_27__data__0__anchor__in;
	assign phi_n26__fork_27__data__0__anchor__out = phi_n26_out1_data;
	assign fork_27_in1_valid = phi_n26__fork_27__valid__0__anchor__in;
	assign phi_n26__fork_27__valid__0__anchor__out = phi_n26_out1_valid;
	assign phi_n26_out1_ready = phi_n26__fork_27__ready__0__anchor__in;
	assign phi_n26__fork_27__ready__0__anchor__out = fork_27_in1_ready;
	assign phi_n27_clk = clk;
	assign phi_n27_rst = rst;
	assign fork_28_in1_data = phi_n27__fork_28__data__0__anchor__in;
	assign phi_n27__fork_28__data__0__anchor__out = phi_n27_out1_data;
	assign fork_28_in1_valid = phi_n27__fork_28__valid__0__anchor__in;
	assign phi_n27__fork_28__valid__0__anchor__out = phi_n27_out1_valid;
	assign phi_n27_out1_ready = phi_n27__fork_28__ready__0__anchor__in;
	assign phi_n27__fork_28__ready__0__anchor__out = fork_28_in1_ready;
	assign fork_0_clk = clk;
	assign fork_0_rst = rst;
	assign add_5_in2_data = fork_0__add_5__data__0__anchor__in;
	assign fork_0__add_5__data__0__anchor__out = fork_0_out1_data;
	assign add_5_in2_valid = fork_0__add_5__valid__0__anchor__in;
	assign fork_0__add_5__valid__0__anchor__out = fork_0_out1_valid;
	assign fork_0_out1_ready = fork_0__add_5__ready__0__anchor__in;
	assign fork_0__add_5__ready__0__anchor__out = add_5_in2_ready;
	assign add_26_in2_data = fork_0__add_26__data__0__anchor__in;
	assign fork_0__add_26__data__0__anchor__out = fork_0_out2_data;
	assign add_26_in2_valid = fork_0__add_26__valid__0__anchor__in;
	assign fork_0__add_26__valid__0__anchor__out = fork_0_out2_valid;
	assign fork_0_out2_ready = fork_0__add_26__ready__0__anchor__in;
	assign fork_0__add_26__ready__0__anchor__out = add_26_in2_ready;
	assign add_29_in1_data = fork_0__add_29__data__0__anchor__in;
	assign fork_0__add_29__data__0__anchor__out = fork_0_out3_data;
	assign add_29_in1_valid = fork_0__add_29__valid__0__anchor__in;
	assign fork_0__add_29__valid__0__anchor__out = fork_0_out3_valid;
	assign fork_0_out3_ready = fork_0__add_29__ready__0__anchor__in;
	assign fork_0__add_29__ready__0__anchor__out = add_29_in1_ready;
	assign load_14_in2_data = fork_0__load_14__data__0__anchor__in;
	assign fork_0__load_14__data__0__anchor__out = fork_0_out4_data;
	assign load_14_in2_valid = fork_0__load_14__valid__0__anchor__in;
	assign fork_0__load_14__valid__0__anchor__out = fork_0_out4_valid;
	assign fork_0_out4_ready = fork_0__load_14__ready__0__anchor__in;
	assign fork_0__load_14__ready__0__anchor__out = load_14_in2_ready;
	assign load_22_in2_data = fork_0__load_22__data__0__anchor__in;
	assign fork_0__load_22__data__0__anchor__out = fork_0_out5_data;
	assign load_22_in2_valid = fork_0__load_22__valid__0__anchor__in;
	assign fork_0__load_22__valid__0__anchor__out = fork_0_out5_valid;
	assign fork_0_out5_ready = fork_0__load_22__ready__0__anchor__in;
	assign fork_0__load_22__ready__0__anchor__out = load_22_in2_ready;
	assign fork_1_clk = clk;
	assign fork_1_rst = rst;
	assign icmp_30_in1_data = fork_1__icmp_30__data__0__anchor__in;
	assign fork_1__icmp_30__data__0__anchor__out = fork_1_out1_data;
	assign icmp_30_in1_valid = fork_1__icmp_30__valid__0__anchor__in;
	assign fork_1__icmp_30__valid__0__anchor__out = fork_1_out1_valid;
	assign fork_1_out1_ready = fork_1__icmp_30__ready__0__anchor__in;
	assign fork_1__icmp_30__ready__0__anchor__out = icmp_30_in1_ready;
	assign branch_7_in1_data = fork_1__branch_7__data__0__anchor__in;
	assign fork_1__branch_7__data__0__anchor__out = fork_1_out2_data;
	assign branch_7_in1_valid = fork_1__branch_7__valid__0__anchor__in;
	assign fork_1__branch_7__valid__0__anchor__out = fork_1_out2_valid;
	assign fork_1_out2_ready = fork_1__branch_7__ready__0__anchor__in;
	assign fork_1__branch_7__ready__0__anchor__out = branch_7_in1_ready;
	assign fork_2_clk = clk;
	assign fork_2_rst = rst;
	assign icmp_33_in1_data = fork_2__icmp_33__data__0__anchor__in;
	assign fork_2__icmp_33__data__0__anchor__out = fork_2_out1_data;
	assign icmp_33_in1_valid = fork_2__icmp_33__valid__0__anchor__in;
	assign fork_2__icmp_33__valid__0__anchor__out = fork_2_out1_valid;
	assign fork_2_out1_ready = fork_2__icmp_33__ready__0__anchor__in;
	assign fork_2__icmp_33__ready__0__anchor__out = icmp_33_in1_ready;
	assign branch_11_in1_data = fork_2__branch_11__data__0__anchor__in;
	assign fork_2__branch_11__data__0__anchor__out = fork_2_out2_data;
	assign branch_11_in1_valid = fork_2__branch_11__valid__0__anchor__in;
	assign fork_2__branch_11__valid__0__anchor__out = fork_2_out2_valid;
	assign fork_2_out2_ready = fork_2__branch_11__ready__0__anchor__in;
	assign fork_2__branch_11__ready__0__anchor__out = branch_11_in1_ready;
	assign fork_3_clk = clk;
	assign fork_3_rst = rst;
	assign load_39_in2_data = fork_3__load_39__data__0__anchor__in;
	assign fork_3__load_39__data__0__anchor__out = fork_3_out1_data;
	assign load_39_in2_valid = fork_3__load_39__valid__0__anchor__in;
	assign fork_3__load_39__valid__0__anchor__out = fork_3_out1_valid;
	assign fork_3_out1_ready = fork_3__load_39__ready__0__anchor__in;
	assign fork_3__load_39__ready__0__anchor__out = load_39_in2_ready;
	assign branch_21_in1_data = fork_3__branch_21__data__0__anchor__in;
	assign fork_3__branch_21__data__0__anchor__out = fork_3_out2_data;
	assign branch_21_in1_valid = fork_3__branch_21__valid__0__anchor__in;
	assign fork_3__branch_21__valid__0__anchor__out = fork_3_out2_valid;
	assign fork_3_out2_ready = fork_3__branch_21__ready__0__anchor__in;
	assign fork_3__branch_21__ready__0__anchor__out = branch_21_in1_ready;
	assign fork_4_clk = clk;
	assign fork_4_rst = rst;
	assign shl_43_in1_data = fork_4__shl_43__data__0__anchor__in;
	assign fork_4__shl_43__data__0__anchor__out = fork_4_out1_data;
	assign shl_43_in1_valid = fork_4__shl_43__valid__0__anchor__in;
	assign fork_4__shl_43__valid__0__anchor__out = fork_4_out1_valid;
	assign fork_4_out1_ready = fork_4__shl_43__ready__0__anchor__in;
	assign fork_4__shl_43__ready__0__anchor__out = shl_43_in1_ready;
	assign add_54_in1_data = fork_4__add_54__data__0__anchor__in;
	assign fork_4__add_54__data__0__anchor__out = fork_4_out2_data;
	assign add_54_in1_valid = fork_4__add_54__valid__0__anchor__in;
	assign fork_4__add_54__valid__0__anchor__out = fork_4_out2_valid;
	assign fork_4_out2_ready = fork_4__add_54__ready__0__anchor__in;
	assign fork_4__add_54__ready__0__anchor__out = add_54_in1_ready;
	assign load_51_in2_data = fork_4__load_51__data__0__anchor__in;
	assign fork_4__load_51__data__0__anchor__out = fork_4_out3_data;
	assign load_51_in2_valid = fork_4__load_51__valid__0__anchor__in;
	assign fork_4__load_51__valid__0__anchor__out = fork_4_out3_valid;
	assign fork_4_out3_ready = fork_4__load_51__ready__0__anchor__in;
	assign fork_4__load_51__ready__0__anchor__out = load_51_in2_ready;
	assign fork_6_clk = clk;
	assign fork_6_rst = rst;
	assign icmp_55_in1_data = fork_6__icmp_55__data__0__anchor__in;
	assign fork_6__icmp_55__data__0__anchor__out = fork_6_out1_data;
	assign icmp_55_in1_valid = fork_6__icmp_55__valid__0__anchor__in;
	assign fork_6__icmp_55__valid__0__anchor__out = fork_6_out1_valid;
	assign fork_6_out1_ready = fork_6__icmp_55__ready__0__anchor__in;
	assign fork_6__icmp_55__ready__0__anchor__out = icmp_55_in1_ready;
	assign branch_23_in1_data = fork_6__branch_23__data__0__anchor__in;
	assign fork_6__branch_23__data__0__anchor__out = fork_6_out2_data;
	assign branch_23_in1_valid = fork_6__branch_23__valid__0__anchor__in;
	assign fork_6__branch_23__valid__0__anchor__out = fork_6_out2_valid;
	assign fork_6_out2_ready = fork_6__branch_23__ready__0__anchor__in;
	assign fork_6__branch_23__ready__0__anchor__out = branch_23_in1_ready;
	assign fork_7_clk = clk;
	assign fork_7_rst = rst;
	assign icmp_60_in1_data = fork_7__icmp_60__data__0__anchor__in;
	assign fork_7__icmp_60__data__0__anchor__out = fork_7_out1_data;
	assign icmp_60_in1_valid = fork_7__icmp_60__valid__0__anchor__in;
	assign fork_7__icmp_60__valid__0__anchor__out = fork_7_out1_valid;
	assign fork_7_out1_ready = fork_7__icmp_60__ready__0__anchor__in;
	assign fork_7__icmp_60__ready__0__anchor__out = icmp_60_in1_ready;
	assign branch_28_in1_data = fork_7__branch_28__data__0__anchor__in;
	assign fork_7__branch_28__data__0__anchor__out = fork_7_out2_data;
	assign branch_28_in1_valid = fork_7__branch_28__valid__0__anchor__in;
	assign fork_7__branch_28__valid__0__anchor__out = fork_7_out2_valid;
	assign fork_7_out2_ready = fork_7__branch_28__ready__0__anchor__in;
	assign fork_7__branch_28__ready__0__anchor__out = branch_28_in1_ready;
	assign fork_8_clk = clk;
	assign fork_8_rst = rst;
	assign add_73_in1_data = fork_8__add_73__data__0__anchor__in;
	assign fork_8__add_73__data__0__anchor__out = fork_8_out1_data;
	assign add_73_in1_valid = fork_8__add_73__valid__0__anchor__in;
	assign fork_8__add_73__valid__0__anchor__out = fork_8_out1_valid;
	assign fork_8_out1_ready = fork_8__add_73__ready__0__anchor__in;
	assign fork_8__add_73__ready__0__anchor__out = add_73_in1_ready;
	assign load_66_in2_data = fork_8__load_66__data__0__anchor__in;
	assign fork_8__load_66__data__0__anchor__out = fork_8_out2_data;
	assign load_66_in2_valid = fork_8__load_66__valid__0__anchor__in;
	assign fork_8__load_66__valid__0__anchor__out = fork_8_out2_valid;
	assign fork_8_out2_ready = fork_8__load_66__ready__0__anchor__in;
	assign fork_8__load_66__ready__0__anchor__out = load_66_in2_ready;
	assign load_69_in2_data = fork_8__load_69__data__0__anchor__in;
	assign fork_8__load_69__data__0__anchor__out = fork_8_out3_data;
	assign load_69_in2_valid = fork_8__load_69__valid__0__anchor__in;
	assign fork_8__load_69__valid__0__anchor__out = fork_8_out3_valid;
	assign fork_8_out3_ready = fork_8__load_69__ready__0__anchor__in;
	assign fork_8__load_69__ready__0__anchor__out = load_69_in2_ready;
	assign store_2_in2_data = fork_8__store_2__data__0__anchor__in;
	assign fork_8__store_2__data__0__anchor__out = fork_8_out4_data;
	assign store_2_in2_valid = fork_8__store_2__valid__0__anchor__in;
	assign fork_8__store_2__valid__0__anchor__out = fork_8_out4_valid;
	assign fork_8_out4_ready = fork_8__store_2__ready__0__anchor__in;
	assign fork_8__store_2__ready__0__anchor__out = store_2_in2_ready;
	assign fork_9_clk = clk;
	assign fork_9_rst = rst;
	assign icmp_74_in1_data = fork_9__icmp_74__data__0__anchor__in;
	assign fork_9__icmp_74__data__0__anchor__out = fork_9_out1_data;
	assign icmp_74_in1_valid = fork_9__icmp_74__valid__0__anchor__in;
	assign fork_9__icmp_74__valid__0__anchor__out = fork_9_out1_valid;
	assign fork_9_out1_ready = fork_9__icmp_74__ready__0__anchor__in;
	assign fork_9__icmp_74__ready__0__anchor__out = icmp_74_in1_ready;
	assign branch_32_in1_data = fork_9__branch_32__data__0__anchor__in;
	assign fork_9__branch_32__data__0__anchor__out = fork_9_out2_data;
	assign branch_32_in1_valid = fork_9__branch_32__valid__0__anchor__in;
	assign fork_9__branch_32__valid__0__anchor__out = fork_9_out2_valid;
	assign fork_9_out2_ready = fork_9__branch_32__ready__0__anchor__in;
	assign fork_9__branch_32__ready__0__anchor__out = branch_32_in1_ready;
	assign fork_10_clk = clk;
	assign fork_10_rst = rst;
	assign load_80_in2_data = fork_10__load_80__data__0__anchor__in;
	assign fork_10__load_80__data__0__anchor__out = fork_10_out1_data;
	assign load_80_in2_valid = fork_10__load_80__valid__0__anchor__in;
	assign fork_10__load_80__valid__0__anchor__out = fork_10_out1_valid;
	assign fork_10_out1_ready = fork_10__load_80__ready__0__anchor__in;
	assign fork_10__load_80__ready__0__anchor__out = load_80_in2_ready;
	assign branch_39_in1_data = fork_10__branch_39__data__0__anchor__in;
	assign fork_10__branch_39__data__0__anchor__out = fork_10_out2_data;
	assign branch_39_in1_valid = fork_10__branch_39__valid__0__anchor__in;
	assign fork_10__branch_39__valid__0__anchor__out = fork_10_out2_valid;
	assign fork_10_out2_ready = fork_10__branch_39__ready__0__anchor__in;
	assign fork_10__branch_39__ready__0__anchor__out = branch_39_in1_ready;
	assign fork_11_clk = clk;
	assign fork_11_rst = rst;
	assign add_85_in2_data = fork_11__add_85__data__0__anchor__in;
	assign fork_11__add_85__data__0__anchor__out = fork_11_out1_data;
	assign add_85_in2_valid = fork_11__add_85__valid__0__anchor__in;
	assign fork_11__add_85__valid__0__anchor__out = fork_11_out1_valid;
	assign fork_11_out1_ready = fork_11__add_85__ready__0__anchor__in;
	assign fork_11__add_85__ready__0__anchor__out = add_85_in2_ready;
	assign add_95_in1_data = fork_11__add_95__data__0__anchor__in;
	assign fork_11__add_95__data__0__anchor__out = fork_11_out2_data;
	assign add_95_in1_valid = fork_11__add_95__valid__0__anchor__in;
	assign fork_11__add_95__valid__0__anchor__out = fork_11_out2_valid;
	assign fork_11_out2_ready = fork_11__add_95__ready__0__anchor__in;
	assign fork_11__add_95__ready__0__anchor__out = add_95_in1_ready;
	assign load_92_in2_data = fork_11__load_92__data__0__anchor__in;
	assign fork_11__load_92__data__0__anchor__out = fork_11_out3_data;
	assign load_92_in2_valid = fork_11__load_92__valid__0__anchor__in;
	assign fork_11__load_92__valid__0__anchor__out = fork_11_out3_valid;
	assign fork_11_out3_ready = fork_11__load_92__ready__0__anchor__in;
	assign fork_11__load_92__ready__0__anchor__out = load_92_in2_ready;
	assign fork_13_clk = clk;
	assign fork_13_rst = rst;
	assign icmp_96_in1_data = fork_13__icmp_96__data__0__anchor__in;
	assign fork_13__icmp_96__data__0__anchor__out = fork_13_out1_data;
	assign icmp_96_in1_valid = fork_13__icmp_96__valid__0__anchor__in;
	assign fork_13__icmp_96__valid__0__anchor__out = fork_13_out1_valid;
	assign fork_13_out1_ready = fork_13__icmp_96__ready__0__anchor__in;
	assign fork_13__icmp_96__ready__0__anchor__out = icmp_96_in1_ready;
	assign branch_41_in1_data = fork_13__branch_41__data__0__anchor__in;
	assign fork_13__branch_41__data__0__anchor__out = fork_13_out2_data;
	assign branch_41_in1_valid = fork_13__branch_41__valid__0__anchor__in;
	assign fork_13__branch_41__valid__0__anchor__out = fork_13_out2_valid;
	assign fork_13_out2_ready = fork_13__branch_41__ready__0__anchor__in;
	assign fork_13__branch_41__ready__0__anchor__out = branch_41_in1_ready;
	assign fork_14_clk = clk;
	assign fork_14_rst = rst;
	assign icmp_101_in1_data = fork_14__icmp_101__data__0__anchor__in;
	assign fork_14__icmp_101__data__0__anchor__out = fork_14_out1_data;
	assign icmp_101_in1_valid = fork_14__icmp_101__valid__0__anchor__in;
	assign fork_14__icmp_101__valid__0__anchor__out = fork_14_out1_valid;
	assign fork_14_out1_ready = fork_14__icmp_101__ready__0__anchor__in;
	assign fork_14__icmp_101__ready__0__anchor__out = icmp_101_in1_ready;
	assign branch_45_in1_data = fork_14__branch_45__data__0__anchor__in;
	assign fork_14__branch_45__data__0__anchor__out = fork_14_out2_data;
	assign branch_45_in1_valid = fork_14__branch_45__valid__0__anchor__in;
	assign fork_14__branch_45__valid__0__anchor__out = fork_14_out2_valid;
	assign fork_14_out2_ready = fork_14__branch_45__ready__0__anchor__in;
	assign fork_14__branch_45__ready__0__anchor__out = branch_45_in1_ready;
	assign fork_17_clk = clk;
	assign fork_17_rst = rst;
	assign shl_4_in1_data = fork_17__shl_4__data__0__anchor__in;
	assign fork_17__shl_4__data__0__anchor__out = fork_17_out1_data;
	assign shl_4_in1_valid = fork_17__shl_4__valid__0__anchor__in;
	assign fork_17__shl_4__valid__0__anchor__out = fork_17_out1_valid;
	assign fork_17_out1_ready = fork_17__shl_4__ready__0__anchor__in;
	assign fork_17__shl_4__ready__0__anchor__out = shl_4_in1_ready;
	assign load_11_in2_data = fork_17__load_11__data__0__anchor__in;
	assign fork_17__load_11__data__0__anchor__out = fork_17_out2_data;
	assign load_11_in2_valid = fork_17__load_11__valid__0__anchor__in;
	assign fork_17__load_11__valid__0__anchor__out = fork_17_out2_valid;
	assign fork_17_out2_ready = fork_17__load_11__ready__0__anchor__in;
	assign fork_17__load_11__ready__0__anchor__out = load_11_in2_ready;
	assign load_19_in2_data = fork_17__load_19__data__0__anchor__in;
	assign fork_17__load_19__data__0__anchor__out = fork_17_out3_data;
	assign load_19_in2_valid = fork_17__load_19__valid__0__anchor__in;
	assign fork_17__load_19__valid__0__anchor__out = fork_17_out3_valid;
	assign fork_17_out3_ready = fork_17__load_19__ready__0__anchor__in;
	assign fork_17__load_19__ready__0__anchor__out = load_19_in2_ready;
	assign shl_25_in1_data = fork_17__shl_25__data__0__anchor__in;
	assign fork_17__shl_25__data__0__anchor__out = fork_17_out4_data;
	assign shl_25_in1_valid = fork_17__shl_25__valid__0__anchor__in;
	assign fork_17__shl_25__valid__0__anchor__out = fork_17_out4_valid;
	assign fork_17_out4_ready = fork_17__shl_25__ready__0__anchor__in;
	assign fork_17__shl_25__ready__0__anchor__out = shl_25_in1_ready;
	assign branch_8_in1_data = fork_17__branch_8__data__0__anchor__in;
	assign fork_17__branch_8__data__0__anchor__out = fork_17_out5_data;
	assign branch_8_in1_valid = fork_17__branch_8__valid__0__anchor__in;
	assign fork_17__branch_8__valid__0__anchor__out = fork_17_out5_valid;
	assign fork_17_out5_ready = fork_17__branch_8__ready__0__anchor__in;
	assign fork_17__branch_8__ready__0__anchor__out = branch_8_in1_ready;
	assign fork_20_clk = clk;
	assign fork_20_rst = rst;
	assign store_1_in2_data = fork_20__store_1__data__0__anchor__in;
	assign fork_20__store_1__data__0__anchor__out = fork_20_out1_data;
	assign store_1_in2_valid = fork_20__store_1__valid__0__anchor__in;
	assign fork_20__store_1__valid__0__anchor__out = fork_20_out1_valid;
	assign fork_20_out1_ready = fork_20__store_1__ready__0__anchor__in;
	assign fork_20__store_1__ready__0__anchor__out = store_1_in2_ready;
	assign add_59_in1_data = fork_20__add_59__data__0__anchor__in;
	assign fork_20__add_59__data__0__anchor__out = fork_20_out2_data;
	assign add_59_in1_valid = fork_20__add_59__valid__0__anchor__in;
	assign fork_20__add_59__valid__0__anchor__out = fork_20_out2_valid;
	assign fork_20_out2_ready = fork_20__add_59__ready__0__anchor__in;
	assign fork_20__add_59__ready__0__anchor__out = add_59_in1_ready;
	assign fork_22_clk = clk;
	assign fork_22_rst = rst;
	assign add_44_in2_data = fork_22__add_44__data__0__anchor__in;
	assign fork_22__add_44__data__0__anchor__out = fork_22_out1_data;
	assign add_44_in2_valid = fork_22__add_44__valid__0__anchor__in;
	assign fork_22__add_44__valid__0__anchor__out = fork_22_out1_valid;
	assign fork_22_out1_ready = fork_22__add_44__ready__0__anchor__in;
	assign fork_22__add_44__ready__0__anchor__out = add_44_in2_ready;
	assign branch_24_in1_data = fork_22__branch_24__data__0__anchor__in;
	assign fork_22__branch_24__data__0__anchor__out = fork_22_out2_data;
	assign branch_24_in1_valid = fork_22__branch_24__valid__0__anchor__in;
	assign fork_22__branch_24__valid__0__anchor__out = fork_22_out2_valid;
	assign fork_22_out2_ready = fork_22__branch_24__ready__0__anchor__in;
	assign fork_22__branch_24__ready__0__anchor__out = branch_24_in1_ready;
	assign fork_23_clk = clk;
	assign fork_23_rst = rst;
	assign mul_48_in2_data = fork_23__mul_48__data__0__anchor__in;
	assign fork_23__mul_48__data__0__anchor__out = fork_23_out1_data;
	assign mul_48_in2_valid = fork_23__mul_48__valid__0__anchor__in;
	assign fork_23__mul_48__valid__0__anchor__out = fork_23_out1_valid;
	assign fork_23_out1_ready = fork_23__mul_48__ready__0__anchor__in;
	assign fork_23__mul_48__ready__0__anchor__out = mul_48_in2_ready;
	assign branch_25_in1_data = fork_23__branch_25__data__0__anchor__in;
	assign fork_23__branch_25__data__0__anchor__out = fork_23_out2_data;
	assign branch_25_in1_valid = fork_23__branch_25__valid__0__anchor__in;
	assign fork_23__branch_25__valid__0__anchor__out = fork_23_out2_valid;
	assign fork_23_out2_ready = fork_23__branch_25__ready__0__anchor__in;
	assign fork_23__branch_25__ready__0__anchor__out = branch_25_in1_ready;
	assign fork_26_clk = clk;
	assign fork_26_rst = rst;
	assign store_3_in2_data = fork_26__store_3__data__0__anchor__in;
	assign fork_26__store_3__data__0__anchor__out = fork_26_out1_data;
	assign store_3_in2_valid = fork_26__store_3__valid__0__anchor__in;
	assign fork_26__store_3__valid__0__anchor__out = fork_26_out1_valid;
	assign fork_26_out1_ready = fork_26__store_3__ready__0__anchor__in;
	assign fork_26__store_3__ready__0__anchor__out = store_3_in2_ready;
	assign add_100_in1_data = fork_26__add_100__data__0__anchor__in;
	assign fork_26__add_100__data__0__anchor__out = fork_26_out2_data;
	assign add_100_in1_valid = fork_26__add_100__valid__0__anchor__in;
	assign fork_26__add_100__valid__0__anchor__out = fork_26_out2_valid;
	assign fork_26_out2_ready = fork_26__add_100__ready__0__anchor__in;
	assign fork_26__add_100__ready__0__anchor__out = add_100_in1_ready;
	assign fork_27_clk = clk;
	assign fork_27_rst = rst;
	assign shl_84_in1_data = fork_27__shl_84__data__0__anchor__in;
	assign fork_27__shl_84__data__0__anchor__out = fork_27_out1_data;
	assign shl_84_in1_valid = fork_27__shl_84__valid__0__anchor__in;
	assign fork_27__shl_84__valid__0__anchor__out = fork_27_out1_valid;
	assign fork_27_out1_ready = fork_27__shl_84__ready__0__anchor__in;
	assign fork_27__shl_84__ready__0__anchor__out = shl_84_in1_ready;
	assign branch_42_in1_data = fork_27__branch_42__data__0__anchor__in;
	assign fork_27__branch_42__data__0__anchor__out = fork_27_out2_data;
	assign branch_42_in1_valid = fork_27__branch_42__valid__0__anchor__in;
	assign fork_27__branch_42__valid__0__anchor__out = fork_27_out2_valid;
	assign fork_27_out2_ready = fork_27__branch_42__ready__0__anchor__in;
	assign fork_27__branch_42__ready__0__anchor__out = branch_42_in1_ready;
	assign fork_28_clk = clk;
	assign fork_28_rst = rst;
	assign mul_89_in2_data = fork_28__mul_89__data__0__anchor__in;
	assign fork_28__mul_89__data__0__anchor__out = fork_28_out1_data;
	assign mul_89_in2_valid = fork_28__mul_89__valid__0__anchor__in;
	assign fork_28__mul_89__valid__0__anchor__out = fork_28_out1_valid;
	assign fork_28_out1_ready = fork_28__mul_89__ready__0__anchor__in;
	assign fork_28__mul_89__ready__0__anchor__out = mul_89_in2_ready;
	assign branch_43_in1_data = fork_28__branch_43__data__0__anchor__in;
	assign fork_28__branch_43__data__0__anchor__out = fork_28_out2_data;
	assign branch_43_in1_valid = fork_28__branch_43__valid__0__anchor__in;
	assign fork_28__branch_43__valid__0__anchor__out = fork_28_out2_valid;
	assign fork_28_out2_ready = fork_28__branch_43__ready__0__anchor__in;
	assign fork_28__branch_43__ready__0__anchor__out = branch_43_in1_ready;
	assign branch_0_clk = clk;
	assign branch_0_rst = rst;
	assign phi_1_in2_data = branch_0__phi_1__data__0__anchor__in;
	assign branch_0__phi_1__data__0__anchor__out = branch_0_out1_data;
	assign phi_1_in2_valid = branch_0__phi_1__valid__0__anchor__in;
	assign branch_0__phi_1__valid__0__anchor__out = branch_0_out1_valid;
	assign branch_0_out1_ready = branch_0__phi_1__ready__0__anchor__in;
	assign branch_0__phi_1__ready__0__anchor__out = phi_1_in2_ready;
	assign sink_0_in1_data = branch_0__sink_0__data__0__anchor__in;
	assign branch_0__sink_0__data__0__anchor__out = branch_0_out2_data;
	assign sink_0_in1_valid = branch_0__sink_0__valid__0__anchor__in;
	assign branch_0__sink_0__valid__0__anchor__out = branch_0_out2_valid;
	assign branch_0_out2_ready = branch_0__sink_0__ready__0__anchor__in;
	assign branch_0__sink_0__ready__0__anchor__out = sink_0_in1_ready;
	assign branch_1_clk = clk;
	assign branch_1_rst = rst;
	assign phi_n0_in1_data = branch_1__phi_n0__data__0__anchor__in;
	assign branch_1__phi_n0__data__0__anchor__out = branch_1_out1_data;
	assign phi_n0_in1_valid = branch_1__phi_n0__valid__0__anchor__in;
	assign branch_1__phi_n0__valid__0__anchor__out = branch_1_out1_valid;
	assign branch_1_out1_ready = branch_1__phi_n0__ready__0__anchor__in;
	assign branch_1__phi_n0__ready__0__anchor__out = phi_n0_in1_ready;
	assign sink_1_in1_data = branch_1__sink_1__data__0__anchor__in;
	assign branch_1__sink_1__data__0__anchor__out = branch_1_out2_data;
	assign sink_1_in1_valid = branch_1__sink_1__valid__0__anchor__in;
	assign branch_1__sink_1__valid__0__anchor__out = branch_1_out2_valid;
	assign branch_1_out2_ready = branch_1__sink_1__ready__0__anchor__in;
	assign branch_1__sink_1__ready__0__anchor__out = sink_1_in1_ready;
	assign branch_2_clk = clk;
	assign branch_2_rst = rst;
	assign phi_n1_in1_data = branch_2__phi_n1__data__0__anchor__in;
	assign branch_2__phi_n1__data__0__anchor__out = branch_2_out1_data;
	assign phi_n1_in1_valid = branch_2__phi_n1__valid__0__anchor__in;
	assign branch_2__phi_n1__valid__0__anchor__out = branch_2_out1_valid;
	assign branch_2_out1_ready = branch_2__phi_n1__ready__0__anchor__in;
	assign branch_2__phi_n1__ready__0__anchor__out = phi_n1_in1_ready;
	assign sink_2_in1_data = branch_2__sink_2__data__0__anchor__in;
	assign branch_2__sink_2__data__0__anchor__out = branch_2_out2_data;
	assign sink_2_in1_valid = branch_2__sink_2__valid__0__anchor__in;
	assign branch_2__sink_2__valid__0__anchor__out = branch_2_out2_valid;
	assign branch_2_out2_ready = branch_2__sink_2__ready__0__anchor__in;
	assign branch_2__sink_2__ready__0__anchor__out = sink_2_in1_ready;
	assign fork_29_clk = clk;
	assign fork_29_rst = rst;
	assign branch_2_in2_data = fork_29__branch_2__data__0__anchor__in;
	assign fork_29__branch_2__data__0__anchor__out = fork_29_out1_data;
	assign branch_2_in2_valid = fork_29__branch_2__valid__0__anchor__in;
	assign fork_29__branch_2__valid__0__anchor__out = fork_29_out1_valid;
	assign fork_29_out1_ready = fork_29__branch_2__ready__0__anchor__in;
	assign fork_29__branch_2__ready__0__anchor__out = branch_2_in2_ready;
	assign branch_1_in2_data = fork_29__branch_1__data__0__anchor__in;
	assign fork_29__branch_1__data__0__anchor__out = fork_29_out2_data;
	assign branch_1_in2_valid = fork_29__branch_1__valid__0__anchor__in;
	assign fork_29__branch_1__valid__0__anchor__out = fork_29_out2_valid;
	assign fork_29_out2_ready = fork_29__branch_1__ready__0__anchor__in;
	assign fork_29__branch_1__ready__0__anchor__out = branch_1_in2_ready;
	assign branch_0_in2_data = fork_29__branch_0__data__0__anchor__in;
	assign fork_29__branch_0__data__0__anchor__out = fork_29_out3_data;
	assign branch_0_in2_valid = fork_29__branch_0__valid__0__anchor__in;
	assign fork_29__branch_0__valid__0__anchor__out = fork_29_out3_valid;
	assign fork_29_out3_ready = fork_29__branch_0__ready__0__anchor__in;
	assign fork_29__branch_0__ready__0__anchor__out = branch_0_in2_ready;
	assign branchC_46_in2_data = fork_29__branchC_46__data__0__anchor__in;
	assign fork_29__branchC_46__data__0__anchor__out = fork_29_out4_data;
	assign branchC_46_in2_valid = fork_29__branchC_46__valid__0__anchor__in;
	assign fork_29__branchC_46__valid__0__anchor__out = fork_29_out4_valid;
	assign fork_29_out4_ready = fork_29__branchC_46__ready__0__anchor__in;
	assign fork_29__branchC_46__ready__0__anchor__out = branchC_46_in2_ready;
	assign branch_3_clk = clk;
	assign branch_3_rst = rst;
	assign phi_3_in2_data = branch_3__phi_3__data__0__anchor__in;
	assign branch_3__phi_3__data__0__anchor__out = branch_3_out1_data;
	assign phi_3_in2_valid = branch_3__phi_3__valid__0__anchor__in;
	assign branch_3__phi_3__valid__0__anchor__out = branch_3_out1_valid;
	assign branch_3_out1_ready = branch_3__phi_3__ready__0__anchor__in;
	assign branch_3__phi_3__ready__0__anchor__out = phi_3_in2_ready;
	assign sink_3_in1_data = branch_3__sink_3__data__0__anchor__in;
	assign branch_3__sink_3__data__0__anchor__out = branch_3_out2_data;
	assign sink_3_in1_valid = branch_3__sink_3__valid__0__anchor__in;
	assign branch_3__sink_3__valid__0__anchor__out = branch_3_out2_valid;
	assign branch_3_out2_ready = branch_3__sink_3__ready__0__anchor__in;
	assign branch_3__sink_3__ready__0__anchor__out = sink_3_in1_ready;
	assign branch_4_clk = clk;
	assign branch_4_rst = rst;
	assign phi_n5_in1_data = branch_4__phi_n5__data__0__anchor__in;
	assign branch_4__phi_n5__data__0__anchor__out = branch_4_out1_data;
	assign phi_n5_in1_valid = branch_4__phi_n5__valid__0__anchor__in;
	assign branch_4__phi_n5__valid__0__anchor__out = branch_4_out1_valid;
	assign branch_4_out1_ready = branch_4__phi_n5__ready__0__anchor__in;
	assign branch_4__phi_n5__ready__0__anchor__out = phi_n5_in1_ready;
	assign sink_4_in1_data = branch_4__sink_4__data__0__anchor__in;
	assign branch_4__sink_4__data__0__anchor__out = branch_4_out2_data;
	assign sink_4_in1_valid = branch_4__sink_4__valid__0__anchor__in;
	assign branch_4__sink_4__valid__0__anchor__out = branch_4_out2_valid;
	assign branch_4_out2_ready = branch_4__sink_4__ready__0__anchor__in;
	assign branch_4__sink_4__ready__0__anchor__out = sink_4_in1_ready;
	assign branch_5_clk = clk;
	assign branch_5_rst = rst;
	assign phi_n6_in1_data = branch_5__phi_n6__data__0__anchor__in;
	assign branch_5__phi_n6__data__0__anchor__out = branch_5_out1_data;
	assign phi_n6_in1_valid = branch_5__phi_n6__valid__0__anchor__in;
	assign branch_5__phi_n6__valid__0__anchor__out = branch_5_out1_valid;
	assign branch_5_out1_ready = branch_5__phi_n6__ready__0__anchor__in;
	assign branch_5__phi_n6__ready__0__anchor__out = phi_n6_in1_ready;
	assign sink_5_in1_data = branch_5__sink_5__data__0__anchor__in;
	assign branch_5__sink_5__data__0__anchor__out = branch_5_out2_data;
	assign sink_5_in1_valid = branch_5__sink_5__valid__0__anchor__in;
	assign branch_5__sink_5__valid__0__anchor__out = branch_5_out2_valid;
	assign branch_5_out2_ready = branch_5__sink_5__ready__0__anchor__in;
	assign branch_5__sink_5__ready__0__anchor__out = sink_5_in1_ready;
	assign branch_6_clk = clk;
	assign branch_6_rst = rst;
	assign phi_n7_in1_data = branch_6__phi_n7__data__0__anchor__in;
	assign branch_6__phi_n7__data__0__anchor__out = branch_6_out1_data;
	assign phi_n7_in1_valid = branch_6__phi_n7__valid__0__anchor__in;
	assign branch_6__phi_n7__valid__0__anchor__out = branch_6_out1_valid;
	assign branch_6_out1_ready = branch_6__phi_n7__ready__0__anchor__in;
	assign branch_6__phi_n7__ready__0__anchor__out = phi_n7_in1_ready;
	assign sink_6_in1_data = branch_6__sink_6__data__0__anchor__in;
	assign branch_6__sink_6__data__0__anchor__out = branch_6_out2_data;
	assign sink_6_in1_valid = branch_6__sink_6__valid__0__anchor__in;
	assign branch_6__sink_6__valid__0__anchor__out = branch_6_out2_valid;
	assign branch_6_out2_ready = branch_6__sink_6__ready__0__anchor__in;
	assign branch_6__sink_6__ready__0__anchor__out = sink_6_in1_ready;
	assign fork_30_clk = clk;
	assign fork_30_rst = rst;
	assign branch_6_in2_data = fork_30__branch_6__data__0__anchor__in;
	assign fork_30__branch_6__data__0__anchor__out = fork_30_out1_data;
	assign branch_6_in2_valid = fork_30__branch_6__valid__0__anchor__in;
	assign fork_30__branch_6__valid__0__anchor__out = fork_30_out1_valid;
	assign fork_30_out1_ready = fork_30__branch_6__ready__0__anchor__in;
	assign fork_30__branch_6__ready__0__anchor__out = branch_6_in2_ready;
	assign branch_5_in2_data = fork_30__branch_5__data__0__anchor__in;
	assign fork_30__branch_5__data__0__anchor__out = fork_30_out2_data;
	assign branch_5_in2_valid = fork_30__branch_5__valid__0__anchor__in;
	assign fork_30__branch_5__valid__0__anchor__out = fork_30_out2_valid;
	assign fork_30_out2_ready = fork_30__branch_5__ready__0__anchor__in;
	assign fork_30__branch_5__ready__0__anchor__out = branch_5_in2_ready;
	assign branch_4_in2_data = fork_30__branch_4__data__0__anchor__in;
	assign fork_30__branch_4__data__0__anchor__out = fork_30_out3_data;
	assign branch_4_in2_valid = fork_30__branch_4__valid__0__anchor__in;
	assign fork_30__branch_4__valid__0__anchor__out = fork_30_out3_valid;
	assign fork_30_out3_ready = fork_30__branch_4__ready__0__anchor__in;
	assign fork_30__branch_4__ready__0__anchor__out = branch_4_in2_ready;
	assign branch_3_in2_data = fork_30__branch_3__data__0__anchor__in;
	assign fork_30__branch_3__data__0__anchor__out = fork_30_out4_data;
	assign branch_3_in2_valid = fork_30__branch_3__valid__0__anchor__in;
	assign fork_30__branch_3__valid__0__anchor__out = fork_30_out4_valid;
	assign fork_30_out4_ready = fork_30__branch_3__ready__0__anchor__in;
	assign fork_30__branch_3__ready__0__anchor__out = branch_3_in2_ready;
	assign branchC_47_in2_data = fork_30__branchC_47__data__0__anchor__in;
	assign fork_30__branchC_47__data__0__anchor__out = fork_30_out5_data;
	assign branchC_47_in2_valid = fork_30__branchC_47__valid__0__anchor__in;
	assign fork_30__branchC_47__valid__0__anchor__out = fork_30_out5_valid;
	assign fork_30_out5_ready = fork_30__branchC_47__ready__0__anchor__in;
	assign fork_30__branchC_47__ready__0__anchor__out = branchC_47_in2_ready;
	assign branch_7_clk = clk;
	assign branch_7_rst = rst;
	assign Buffer_25_in1_data = branch_7__Buffer_25__data__0__anchor__in;
	assign branch_7__Buffer_25__data__0__anchor__out = branch_7_out1_data;
	assign Buffer_25_in1_valid = branch_7__Buffer_25__valid__0__anchor__in;
	assign branch_7__Buffer_25__valid__0__anchor__out = branch_7_out1_valid;
	assign branch_7_out1_ready = branch_7__Buffer_25__ready__0__anchor__in;
	assign branch_7__Buffer_25__ready__0__anchor__out = Buffer_25_in1_ready;
	assign sink_7_in1_data = branch_7__sink_7__data__0__anchor__in;
	assign branch_7__sink_7__data__0__anchor__out = branch_7_out2_data;
	assign sink_7_in1_valid = branch_7__sink_7__valid__0__anchor__in;
	assign branch_7__sink_7__valid__0__anchor__out = branch_7_out2_valid;
	assign branch_7_out2_ready = branch_7__sink_7__ready__0__anchor__in;
	assign branch_7__sink_7__ready__0__anchor__out = sink_7_in1_ready;
	assign branch_8_clk = clk;
	assign branch_8_rst = rst;
	assign Buffer_14_in1_data = branch_8__Buffer_14__data__0__anchor__in;
	assign branch_8__Buffer_14__data__0__anchor__out = branch_8_out1_data;
	assign Buffer_14_in1_valid = branch_8__Buffer_14__valid__0__anchor__in;
	assign branch_8__Buffer_14__valid__0__anchor__out = branch_8_out1_valid;
	assign branch_8_out1_ready = branch_8__Buffer_14__ready__0__anchor__in;
	assign branch_8__Buffer_14__ready__0__anchor__out = Buffer_14_in1_ready;
	assign phi_n2_in1_data = branch_8__phi_n2__data__0__anchor__in;
	assign branch_8__phi_n2__data__0__anchor__out = branch_8_out2_data;
	assign phi_n2_in1_valid = branch_8__phi_n2__valid__0__anchor__in;
	assign branch_8__phi_n2__valid__0__anchor__out = branch_8_out2_valid;
	assign branch_8_out2_ready = branch_8__phi_n2__ready__0__anchor__in;
	assign branch_8__phi_n2__ready__0__anchor__out = phi_n2_in1_ready;
	assign branch_9_clk = clk;
	assign branch_9_rst = rst;
	assign Buffer_4_in1_data = branch_9__Buffer_4__data__0__anchor__in;
	assign branch_9__Buffer_4__data__0__anchor__out = branch_9_out1_data;
	assign Buffer_4_in1_valid = branch_9__Buffer_4__valid__0__anchor__in;
	assign branch_9__Buffer_4__valid__0__anchor__out = branch_9_out1_valid;
	assign branch_9_out1_ready = branch_9__Buffer_4__ready__0__anchor__in;
	assign branch_9__Buffer_4__ready__0__anchor__out = Buffer_4_in1_ready;
	assign phi_n3_in1_data = branch_9__phi_n3__data__0__anchor__in;
	assign branch_9__phi_n3__data__0__anchor__out = branch_9_out2_data;
	assign phi_n3_in1_valid = branch_9__phi_n3__valid__0__anchor__in;
	assign branch_9__phi_n3__valid__0__anchor__out = branch_9_out2_valid;
	assign branch_9_out2_ready = branch_9__phi_n3__ready__0__anchor__in;
	assign branch_9__phi_n3__ready__0__anchor__out = phi_n3_in1_ready;
	assign branch_10_clk = clk;
	assign branch_10_rst = rst;
	assign Buffer_5_in1_data = branch_10__Buffer_5__data__0__anchor__in;
	assign branch_10__Buffer_5__data__0__anchor__out = branch_10_out1_data;
	assign Buffer_5_in1_valid = branch_10__Buffer_5__valid__0__anchor__in;
	assign branch_10__Buffer_5__valid__0__anchor__out = branch_10_out1_valid;
	assign branch_10_out1_ready = branch_10__Buffer_5__ready__0__anchor__in;
	assign branch_10__Buffer_5__ready__0__anchor__out = Buffer_5_in1_ready;
	assign phi_n4_in1_data = branch_10__phi_n4__data__0__anchor__in;
	assign branch_10__phi_n4__data__0__anchor__out = branch_10_out2_data;
	assign phi_n4_in1_valid = branch_10__phi_n4__valid__0__anchor__in;
	assign branch_10__phi_n4__valid__0__anchor__out = branch_10_out2_valid;
	assign branch_10_out2_ready = branch_10__phi_n4__ready__0__anchor__in;
	assign branch_10__phi_n4__ready__0__anchor__out = phi_n4_in1_ready;
	assign fork_31_clk = clk;
	assign fork_31_rst = rst;
	assign branch_10_in2_data = fork_31__branch_10__data__0__anchor__in;
	assign fork_31__branch_10__data__0__anchor__out = fork_31_out1_data;
	assign branch_10_in2_valid = fork_31__branch_10__valid__0__anchor__in;
	assign fork_31__branch_10__valid__0__anchor__out = fork_31_out1_valid;
	assign fork_31_out1_ready = fork_31__branch_10__ready__0__anchor__in;
	assign fork_31__branch_10__ready__0__anchor__out = branch_10_in2_ready;
	assign branch_9_in2_data = fork_31__branch_9__data__0__anchor__in;
	assign fork_31__branch_9__data__0__anchor__out = fork_31_out2_data;
	assign branch_9_in2_valid = fork_31__branch_9__valid__0__anchor__in;
	assign fork_31__branch_9__valid__0__anchor__out = fork_31_out2_valid;
	assign fork_31_out2_ready = fork_31__branch_9__ready__0__anchor__in;
	assign fork_31__branch_9__ready__0__anchor__out = branch_9_in2_ready;
	assign branch_8_in2_data = fork_31__branch_8__data__0__anchor__in;
	assign fork_31__branch_8__data__0__anchor__out = fork_31_out3_data;
	assign branch_8_in2_valid = fork_31__branch_8__valid__0__anchor__in;
	assign fork_31__branch_8__valid__0__anchor__out = fork_31_out3_valid;
	assign fork_31_out3_ready = fork_31__branch_8__ready__0__anchor__in;
	assign fork_31__branch_8__ready__0__anchor__out = branch_8_in2_ready;
	assign branch_7_in2_data = fork_31__branch_7__data__0__anchor__in;
	assign fork_31__branch_7__data__0__anchor__out = fork_31_out4_data;
	assign branch_7_in2_valid = fork_31__branch_7__valid__0__anchor__in;
	assign fork_31__branch_7__valid__0__anchor__out = fork_31_out4_valid;
	assign fork_31_out4_ready = fork_31__branch_7__ready__0__anchor__in;
	assign fork_31__branch_7__ready__0__anchor__out = branch_7_in2_ready;
	assign branchC_48_in2_data = fork_31__branchC_48__data__0__anchor__in;
	assign fork_31__branchC_48__data__0__anchor__out = fork_31_out5_data;
	assign branchC_48_in2_valid = fork_31__branchC_48__valid__0__anchor__in;
	assign fork_31__branchC_48__valid__0__anchor__out = fork_31_out5_valid;
	assign fork_31_out5_ready = fork_31__branchC_48__ready__0__anchor__in;
	assign fork_31__branchC_48__ready__0__anchor__out = branchC_48_in2_ready;
	assign branch_11_clk = clk;
	assign branch_11_rst = rst;
	assign Buffer_26_in1_data = branch_11__Buffer_26__data__0__anchor__in;
	assign branch_11__Buffer_26__data__0__anchor__out = branch_11_out1_data;
	assign Buffer_26_in1_valid = branch_11__Buffer_26__valid__0__anchor__in;
	assign branch_11__Buffer_26__valid__0__anchor__out = branch_11_out1_valid;
	assign branch_11_out1_ready = branch_11__Buffer_26__ready__0__anchor__in;
	assign branch_11__Buffer_26__ready__0__anchor__out = Buffer_26_in1_ready;
	assign sink_8_in1_data = branch_11__sink_8__data__0__anchor__in;
	assign branch_11__sink_8__data__0__anchor__out = branch_11_out2_data;
	assign sink_8_in1_valid = branch_11__sink_8__valid__0__anchor__in;
	assign branch_11__sink_8__valid__0__anchor__out = branch_11_out2_valid;
	assign branch_11_out2_ready = branch_11__sink_8__ready__0__anchor__in;
	assign branch_11__sink_8__ready__0__anchor__out = sink_8_in1_ready;
	assign branch_12_clk = clk;
	assign branch_12_rst = rst;
	assign Buffer_1_in1_data = branch_12__Buffer_1__data__0__anchor__in;
	assign branch_12__Buffer_1__data__0__anchor__out = branch_12_out1_data;
	assign Buffer_1_in1_valid = branch_12__Buffer_1__valid__0__anchor__in;
	assign branch_12__Buffer_1__valid__0__anchor__out = branch_12_out1_valid;
	assign branch_12_out1_ready = branch_12__Buffer_1__ready__0__anchor__in;
	assign branch_12__Buffer_1__ready__0__anchor__out = Buffer_1_in1_ready;
	assign phi_n8_in1_data = branch_12__phi_n8__data__0__anchor__in;
	assign branch_12__phi_n8__data__0__anchor__out = branch_12_out2_data;
	assign phi_n8_in1_valid = branch_12__phi_n8__valid__0__anchor__in;
	assign branch_12__phi_n8__valid__0__anchor__out = branch_12_out2_valid;
	assign branch_12_out2_ready = branch_12__phi_n8__ready__0__anchor__in;
	assign branch_12__phi_n8__ready__0__anchor__out = phi_n8_in1_ready;
	assign branch_13_clk = clk;
	assign branch_13_rst = rst;
	assign Buffer_19_in1_data = branch_13__Buffer_19__data__0__anchor__in;
	assign branch_13__Buffer_19__data__0__anchor__out = branch_13_out1_data;
	assign Buffer_19_in1_valid = branch_13__Buffer_19__valid__0__anchor__in;
	assign branch_13__Buffer_19__valid__0__anchor__out = branch_13_out1_valid;
	assign branch_13_out1_ready = branch_13__Buffer_19__ready__0__anchor__in;
	assign branch_13__Buffer_19__ready__0__anchor__out = Buffer_19_in1_ready;
	assign phi_n9_in1_data = branch_13__phi_n9__data__0__anchor__in;
	assign branch_13__phi_n9__data__0__anchor__out = branch_13_out2_data;
	assign phi_n9_in1_valid = branch_13__phi_n9__valid__0__anchor__in;
	assign branch_13__phi_n9__valid__0__anchor__out = branch_13_out2_valid;
	assign branch_13_out2_ready = branch_13__phi_n9__ready__0__anchor__in;
	assign branch_13__phi_n9__ready__0__anchor__out = phi_n9_in1_ready;
	assign fork_32_clk = clk;
	assign fork_32_rst = rst;
	assign branch_13_in2_data = fork_32__branch_13__data__0__anchor__in;
	assign fork_32__branch_13__data__0__anchor__out = fork_32_out1_data;
	assign branch_13_in2_valid = fork_32__branch_13__valid__0__anchor__in;
	assign fork_32__branch_13__valid__0__anchor__out = fork_32_out1_valid;
	assign fork_32_out1_ready = fork_32__branch_13__ready__0__anchor__in;
	assign fork_32__branch_13__ready__0__anchor__out = branch_13_in2_ready;
	assign branch_12_in2_data = fork_32__branch_12__data__0__anchor__in;
	assign fork_32__branch_12__data__0__anchor__out = fork_32_out2_data;
	assign branch_12_in2_valid = fork_32__branch_12__valid__0__anchor__in;
	assign fork_32__branch_12__valid__0__anchor__out = fork_32_out2_valid;
	assign fork_32_out2_ready = fork_32__branch_12__ready__0__anchor__in;
	assign fork_32__branch_12__ready__0__anchor__out = branch_12_in2_ready;
	assign branch_11_in2_data = fork_32__branch_11__data__0__anchor__in;
	assign fork_32__branch_11__data__0__anchor__out = fork_32_out3_data;
	assign branch_11_in2_valid = fork_32__branch_11__valid__0__anchor__in;
	assign fork_32__branch_11__valid__0__anchor__out = fork_32_out3_valid;
	assign fork_32_out3_ready = fork_32__branch_11__ready__0__anchor__in;
	assign fork_32__branch_11__ready__0__anchor__out = branch_11_in2_ready;
	assign branchC_49_in2_data = fork_32__branchC_49__data__0__anchor__in;
	assign fork_32__branchC_49__data__0__anchor__out = fork_32_out4_data;
	assign branchC_49_in2_valid = fork_32__branchC_49__valid__0__anchor__in;
	assign fork_32__branchC_49__valid__0__anchor__out = fork_32_out4_valid;
	assign fork_32_out4_ready = fork_32__branchC_49__ready__0__anchor__in;
	assign fork_32__branchC_49__ready__0__anchor__out = branchC_49_in2_ready;
	assign branch_14_clk = clk;
	assign branch_14_rst = rst;
	assign phi_36_in2_data = branch_14__phi_36__data__0__anchor__in;
	assign branch_14__phi_36__data__0__anchor__out = branch_14_out1_data;
	assign phi_36_in2_valid = branch_14__phi_36__valid__0__anchor__in;
	assign branch_14__phi_36__valid__0__anchor__out = branch_14_out1_valid;
	assign branch_14_out1_ready = branch_14__phi_36__ready__0__anchor__in;
	assign branch_14__phi_36__ready__0__anchor__out = phi_36_in2_ready;
	assign sink_9_in1_data = branch_14__sink_9__data__0__anchor__in;
	assign branch_14__sink_9__data__0__anchor__out = branch_14_out2_data;
	assign sink_9_in1_valid = branch_14__sink_9__valid__0__anchor__in;
	assign branch_14__sink_9__valid__0__anchor__out = branch_14_out2_valid;
	assign branch_14_out2_ready = branch_14__sink_9__ready__0__anchor__in;
	assign branch_14__sink_9__ready__0__anchor__out = sink_9_in1_ready;
	assign branch_15_clk = clk;
	assign branch_15_rst = rst;
	assign phi_n10_in1_data = branch_15__phi_n10__data__0__anchor__in;
	assign branch_15__phi_n10__data__0__anchor__out = branch_15_out1_data;
	assign phi_n10_in1_valid = branch_15__phi_n10__valid__0__anchor__in;
	assign branch_15__phi_n10__valid__0__anchor__out = branch_15_out1_valid;
	assign branch_15_out1_ready = branch_15__phi_n10__ready__0__anchor__in;
	assign branch_15__phi_n10__ready__0__anchor__out = phi_n10_in1_ready;
	assign sink_10_in1_data = branch_15__sink_10__data__0__anchor__in;
	assign branch_15__sink_10__data__0__anchor__out = branch_15_out2_data;
	assign sink_10_in1_valid = branch_15__sink_10__valid__0__anchor__in;
	assign branch_15__sink_10__valid__0__anchor__out = branch_15_out2_valid;
	assign branch_15_out2_ready = branch_15__sink_10__ready__0__anchor__in;
	assign branch_15__sink_10__ready__0__anchor__out = sink_10_in1_ready;
	assign branch_16_clk = clk;
	assign branch_16_rst = rst;
	assign phi_n11_in1_data = branch_16__phi_n11__data__0__anchor__in;
	assign branch_16__phi_n11__data__0__anchor__out = branch_16_out1_data;
	assign phi_n11_in1_valid = branch_16__phi_n11__valid__0__anchor__in;
	assign branch_16__phi_n11__valid__0__anchor__out = branch_16_out1_valid;
	assign branch_16_out1_ready = branch_16__phi_n11__ready__0__anchor__in;
	assign branch_16__phi_n11__ready__0__anchor__out = phi_n11_in1_ready;
	assign sink_11_in1_data = branch_16__sink_11__data__0__anchor__in;
	assign branch_16__sink_11__data__0__anchor__out = branch_16_out2_data;
	assign sink_11_in1_valid = branch_16__sink_11__valid__0__anchor__in;
	assign branch_16__sink_11__valid__0__anchor__out = branch_16_out2_valid;
	assign branch_16_out2_ready = branch_16__sink_11__ready__0__anchor__in;
	assign branch_16__sink_11__ready__0__anchor__out = sink_11_in1_ready;
	assign fork_33_clk = clk;
	assign fork_33_rst = rst;
	assign branch_16_in2_data = fork_33__branch_16__data__0__anchor__in;
	assign fork_33__branch_16__data__0__anchor__out = fork_33_out1_data;
	assign branch_16_in2_valid = fork_33__branch_16__valid__0__anchor__in;
	assign fork_33__branch_16__valid__0__anchor__out = fork_33_out1_valid;
	assign fork_33_out1_ready = fork_33__branch_16__ready__0__anchor__in;
	assign fork_33__branch_16__ready__0__anchor__out = branch_16_in2_ready;
	assign branch_15_in2_data = fork_33__branch_15__data__0__anchor__in;
	assign fork_33__branch_15__data__0__anchor__out = fork_33_out2_data;
	assign branch_15_in2_valid = fork_33__branch_15__valid__0__anchor__in;
	assign fork_33__branch_15__valid__0__anchor__out = fork_33_out2_valid;
	assign fork_33_out2_ready = fork_33__branch_15__ready__0__anchor__in;
	assign fork_33__branch_15__ready__0__anchor__out = branch_15_in2_ready;
	assign branch_14_in2_data = fork_33__branch_14__data__0__anchor__in;
	assign fork_33__branch_14__data__0__anchor__out = fork_33_out3_data;
	assign branch_14_in2_valid = fork_33__branch_14__valid__0__anchor__in;
	assign fork_33__branch_14__valid__0__anchor__out = fork_33_out3_valid;
	assign fork_33_out3_ready = fork_33__branch_14__ready__0__anchor__in;
	assign fork_33__branch_14__ready__0__anchor__out = branch_14_in2_ready;
	assign branchC_50_in2_data = fork_33__branchC_50__data__0__anchor__in;
	assign fork_33__branchC_50__data__0__anchor__out = fork_33_out4_data;
	assign branchC_50_in2_valid = fork_33__branchC_50__valid__0__anchor__in;
	assign fork_33__branchC_50__valid__0__anchor__out = fork_33_out4_valid;
	assign fork_33_out4_ready = fork_33__branchC_50__ready__0__anchor__in;
	assign fork_33__branchC_50__ready__0__anchor__out = branchC_50_in2_ready;
	assign branch_17_clk = clk;
	assign branch_17_rst = rst;
	assign phi_41_in2_data = branch_17__phi_41__data__0__anchor__in;
	assign branch_17__phi_41__data__0__anchor__out = branch_17_out1_data;
	assign phi_41_in2_valid = branch_17__phi_41__valid__0__anchor__in;
	assign branch_17__phi_41__valid__0__anchor__out = branch_17_out1_valid;
	assign branch_17_out1_ready = branch_17__phi_41__ready__0__anchor__in;
	assign branch_17__phi_41__ready__0__anchor__out = phi_41_in2_ready;
	assign sink_12_in1_data = branch_17__sink_12__data__0__anchor__in;
	assign branch_17__sink_12__data__0__anchor__out = branch_17_out2_data;
	assign sink_12_in1_valid = branch_17__sink_12__valid__0__anchor__in;
	assign branch_17__sink_12__valid__0__anchor__out = branch_17_out2_valid;
	assign branch_17_out2_ready = branch_17__sink_12__ready__0__anchor__in;
	assign branch_17__sink_12__ready__0__anchor__out = sink_12_in1_ready;
	assign branch_18_clk = clk;
	assign branch_18_rst = rst;
	assign phi_42_in2_data = branch_18__phi_42__data__0__anchor__in;
	assign branch_18__phi_42__data__0__anchor__out = branch_18_out1_data;
	assign phi_42_in2_valid = branch_18__phi_42__valid__0__anchor__in;
	assign branch_18__phi_42__valid__0__anchor__out = branch_18_out1_valid;
	assign branch_18_out1_ready = branch_18__phi_42__ready__0__anchor__in;
	assign branch_18__phi_42__ready__0__anchor__out = phi_42_in2_ready;
	assign sink_13_in1_data = branch_18__sink_13__data__0__anchor__in;
	assign branch_18__sink_13__data__0__anchor__out = branch_18_out2_data;
	assign sink_13_in1_valid = branch_18__sink_13__valid__0__anchor__in;
	assign branch_18__sink_13__valid__0__anchor__out = branch_18_out2_valid;
	assign branch_18_out2_ready = branch_18__sink_13__ready__0__anchor__in;
	assign branch_18__sink_13__ready__0__anchor__out = sink_13_in1_ready;
	assign branch_19_clk = clk;
	assign branch_19_rst = rst;
	assign phi_n17_in1_data = branch_19__phi_n17__data__0__anchor__in;
	assign branch_19__phi_n17__data__0__anchor__out = branch_19_out1_data;
	assign phi_n17_in1_valid = branch_19__phi_n17__valid__0__anchor__in;
	assign branch_19__phi_n17__valid__0__anchor__out = branch_19_out1_valid;
	assign branch_19_out1_ready = branch_19__phi_n17__ready__0__anchor__in;
	assign branch_19__phi_n17__ready__0__anchor__out = phi_n17_in1_ready;
	assign sink_14_in1_data = branch_19__sink_14__data__0__anchor__in;
	assign branch_19__sink_14__data__0__anchor__out = branch_19_out2_data;
	assign sink_14_in1_valid = branch_19__sink_14__valid__0__anchor__in;
	assign branch_19__sink_14__valid__0__anchor__out = branch_19_out2_valid;
	assign branch_19_out2_ready = branch_19__sink_14__ready__0__anchor__in;
	assign branch_19__sink_14__ready__0__anchor__out = sink_14_in1_ready;
	assign branch_20_clk = clk;
	assign branch_20_rst = rst;
	assign phi_n18_in1_data = branch_20__phi_n18__data__0__anchor__in;
	assign branch_20__phi_n18__data__0__anchor__out = branch_20_out1_data;
	assign phi_n18_in1_valid = branch_20__phi_n18__valid__0__anchor__in;
	assign branch_20__phi_n18__valid__0__anchor__out = branch_20_out1_valid;
	assign branch_20_out1_ready = branch_20__phi_n18__ready__0__anchor__in;
	assign branch_20__phi_n18__ready__0__anchor__out = phi_n18_in1_ready;
	assign sink_15_in1_data = branch_20__sink_15__data__0__anchor__in;
	assign branch_20__sink_15__data__0__anchor__out = branch_20_out2_data;
	assign sink_15_in1_valid = branch_20__sink_15__valid__0__anchor__in;
	assign branch_20__sink_15__valid__0__anchor__out = branch_20_out2_valid;
	assign branch_20_out2_ready = branch_20__sink_15__ready__0__anchor__in;
	assign branch_20__sink_15__ready__0__anchor__out = sink_15_in1_ready;
	assign branch_21_clk = clk;
	assign branch_21_rst = rst;
	assign phi_n16_in1_data = branch_21__phi_n16__data__0__anchor__in;
	assign branch_21__phi_n16__data__0__anchor__out = branch_21_out1_data;
	assign phi_n16_in1_valid = branch_21__phi_n16__valid__0__anchor__in;
	assign branch_21__phi_n16__valid__0__anchor__out = branch_21_out1_valid;
	assign branch_21_out1_ready = branch_21__phi_n16__ready__0__anchor__in;
	assign branch_21__phi_n16__ready__0__anchor__out = phi_n16_in1_ready;
	assign sink_16_in1_data = branch_21__sink_16__data__0__anchor__in;
	assign branch_21__sink_16__data__0__anchor__out = branch_21_out2_data;
	assign sink_16_in1_valid = branch_21__sink_16__valid__0__anchor__in;
	assign branch_21__sink_16__valid__0__anchor__out = branch_21_out2_valid;
	assign branch_21_out2_ready = branch_21__sink_16__ready__0__anchor__in;
	assign branch_21__sink_16__ready__0__anchor__out = sink_16_in1_ready;
	assign fork_34_clk = clk;
	assign fork_34_rst = rst;
	assign branch_21_in2_data = fork_34__branch_21__data__0__anchor__in;
	assign fork_34__branch_21__data__0__anchor__out = fork_34_out1_data;
	assign branch_21_in2_valid = fork_34__branch_21__valid__0__anchor__in;
	assign fork_34__branch_21__valid__0__anchor__out = fork_34_out1_valid;
	assign fork_34_out1_ready = fork_34__branch_21__ready__0__anchor__in;
	assign fork_34__branch_21__ready__0__anchor__out = branch_21_in2_ready;
	assign branch_20_in2_data = fork_34__branch_20__data__0__anchor__in;
	assign fork_34__branch_20__data__0__anchor__out = fork_34_out2_data;
	assign branch_20_in2_valid = fork_34__branch_20__valid__0__anchor__in;
	assign fork_34__branch_20__valid__0__anchor__out = fork_34_out2_valid;
	assign fork_34_out2_ready = fork_34__branch_20__ready__0__anchor__in;
	assign fork_34__branch_20__ready__0__anchor__out = branch_20_in2_ready;
	assign branch_19_in2_data = fork_34__branch_19__data__0__anchor__in;
	assign fork_34__branch_19__data__0__anchor__out = fork_34_out3_data;
	assign branch_19_in2_valid = fork_34__branch_19__valid__0__anchor__in;
	assign fork_34__branch_19__valid__0__anchor__out = fork_34_out3_valid;
	assign fork_34_out3_ready = fork_34__branch_19__ready__0__anchor__in;
	assign fork_34__branch_19__ready__0__anchor__out = branch_19_in2_ready;
	assign branch_18_in2_data = fork_34__branch_18__data__0__anchor__in;
	assign fork_34__branch_18__data__0__anchor__out = fork_34_out4_data;
	assign branch_18_in2_valid = fork_34__branch_18__valid__0__anchor__in;
	assign fork_34__branch_18__valid__0__anchor__out = fork_34_out4_valid;
	assign fork_34_out4_ready = fork_34__branch_18__ready__0__anchor__in;
	assign fork_34__branch_18__ready__0__anchor__out = branch_18_in2_ready;
	assign branch_17_in2_data = fork_34__branch_17__data__0__anchor__in;
	assign fork_34__branch_17__data__0__anchor__out = fork_34_out5_data;
	assign branch_17_in2_valid = fork_34__branch_17__valid__0__anchor__in;
	assign fork_34__branch_17__valid__0__anchor__out = fork_34_out5_valid;
	assign fork_34_out5_ready = fork_34__branch_17__ready__0__anchor__in;
	assign fork_34__branch_17__ready__0__anchor__out = branch_17_in2_ready;
	assign branchC_51_in2_data = fork_34__branchC_51__data__0__anchor__in;
	assign fork_34__branchC_51__data__0__anchor__out = fork_34_out6_data;
	assign branchC_51_in2_valid = fork_34__branchC_51__valid__0__anchor__in;
	assign fork_34__branchC_51__valid__0__anchor__out = fork_34_out6_valid;
	assign fork_34_out6_ready = fork_34__branchC_51__ready__0__anchor__in;
	assign fork_34__branchC_51__ready__0__anchor__out = branchC_51_in2_ready;
	assign branch_22_clk = clk;
	assign branch_22_rst = rst;
	assign Buffer_12_in1_data = branch_22__Buffer_12__data__0__anchor__in;
	assign branch_22__Buffer_12__data__0__anchor__out = branch_22_out1_data;
	assign Buffer_12_in1_valid = branch_22__Buffer_12__valid__0__anchor__in;
	assign branch_22__Buffer_12__valid__0__anchor__out = branch_22_out1_valid;
	assign branch_22_out1_ready = branch_22__Buffer_12__ready__0__anchor__in;
	assign branch_22__Buffer_12__ready__0__anchor__out = Buffer_12_in1_ready;
	assign phi_n12_in1_data = branch_22__phi_n12__data__0__anchor__in;
	assign branch_22__phi_n12__data__0__anchor__out = branch_22_out2_data;
	assign phi_n12_in1_valid = branch_22__phi_n12__valid__0__anchor__in;
	assign branch_22__phi_n12__valid__0__anchor__out = branch_22_out2_valid;
	assign branch_22_out2_ready = branch_22__phi_n12__ready__0__anchor__in;
	assign branch_22__phi_n12__ready__0__anchor__out = phi_n12_in1_ready;
	assign branch_23_clk = clk;
	assign branch_23_rst = rst;
	assign Buffer_3_in1_data = branch_23__Buffer_3__data__0__anchor__in;
	assign branch_23__Buffer_3__data__0__anchor__out = branch_23_out1_data;
	assign Buffer_3_in1_valid = branch_23__Buffer_3__valid__0__anchor__in;
	assign branch_23__Buffer_3__valid__0__anchor__out = branch_23_out1_valid;
	assign branch_23_out1_ready = branch_23__Buffer_3__ready__0__anchor__in;
	assign branch_23__Buffer_3__ready__0__anchor__out = Buffer_3_in1_ready;
	assign sink_17_in1_data = branch_23__sink_17__data__0__anchor__in;
	assign branch_23__sink_17__data__0__anchor__out = branch_23_out2_data;
	assign sink_17_in1_valid = branch_23__sink_17__valid__0__anchor__in;
	assign branch_23__sink_17__valid__0__anchor__out = branch_23_out2_valid;
	assign branch_23_out2_ready = branch_23__sink_17__ready__0__anchor__in;
	assign branch_23__sink_17__ready__0__anchor__out = sink_17_in1_ready;
	assign branch_24_clk = clk;
	assign branch_24_rst = rst;
	assign Buffer_17_in1_data = branch_24__Buffer_17__data__0__anchor__in;
	assign branch_24__Buffer_17__data__0__anchor__out = branch_24_out1_data;
	assign Buffer_17_in1_valid = branch_24__Buffer_17__valid__0__anchor__in;
	assign branch_24__Buffer_17__valid__0__anchor__out = branch_24_out1_valid;
	assign branch_24_out1_ready = branch_24__Buffer_17__ready__0__anchor__in;
	assign branch_24__Buffer_17__ready__0__anchor__out = Buffer_17_in1_ready;
	assign phi_n13_in1_data = branch_24__phi_n13__data__0__anchor__in;
	assign branch_24__phi_n13__data__0__anchor__out = branch_24_out2_data;
	assign phi_n13_in1_valid = branch_24__phi_n13__valid__0__anchor__in;
	assign branch_24__phi_n13__valid__0__anchor__out = branch_24_out2_valid;
	assign branch_24_out2_ready = branch_24__phi_n13__ready__0__anchor__in;
	assign branch_24__phi_n13__ready__0__anchor__out = phi_n13_in1_ready;
	assign branch_25_clk = clk;
	assign branch_25_rst = rst;
	assign Buffer_22_in1_data = branch_25__Buffer_22__data__0__anchor__in;
	assign branch_25__Buffer_22__data__0__anchor__out = branch_25_out1_data;
	assign Buffer_22_in1_valid = branch_25__Buffer_22__valid__0__anchor__in;
	assign branch_25__Buffer_22__valid__0__anchor__out = branch_25_out1_valid;
	assign branch_25_out1_ready = branch_25__Buffer_22__ready__0__anchor__in;
	assign branch_25__Buffer_22__ready__0__anchor__out = Buffer_22_in1_ready;
	assign phi_n14_in1_data = branch_25__phi_n14__data__0__anchor__in;
	assign branch_25__phi_n14__data__0__anchor__out = branch_25_out2_data;
	assign phi_n14_in1_valid = branch_25__phi_n14__valid__0__anchor__in;
	assign branch_25__phi_n14__valid__0__anchor__out = branch_25_out2_valid;
	assign branch_25_out2_ready = branch_25__phi_n14__ready__0__anchor__in;
	assign branch_25__phi_n14__ready__0__anchor__out = phi_n14_in1_ready;
	assign branch_26_clk = clk;
	assign branch_26_rst = rst;
	assign Buffer_18_in1_data = branch_26__Buffer_18__data__0__anchor__in;
	assign branch_26__Buffer_18__data__0__anchor__out = branch_26_out1_data;
	assign Buffer_18_in1_valid = branch_26__Buffer_18__valid__0__anchor__in;
	assign branch_26__Buffer_18__valid__0__anchor__out = branch_26_out1_valid;
	assign branch_26_out1_ready = branch_26__Buffer_18__ready__0__anchor__in;
	assign branch_26__Buffer_18__ready__0__anchor__out = Buffer_18_in1_ready;
	assign phi_n15_in1_data = branch_26__phi_n15__data__0__anchor__in;
	assign branch_26__phi_n15__data__0__anchor__out = branch_26_out2_data;
	assign phi_n15_in1_valid = branch_26__phi_n15__valid__0__anchor__in;
	assign branch_26__phi_n15__valid__0__anchor__out = branch_26_out2_valid;
	assign branch_26_out2_ready = branch_26__phi_n15__ready__0__anchor__in;
	assign branch_26__phi_n15__ready__0__anchor__out = phi_n15_in1_ready;
	assign fork_35_clk = clk;
	assign fork_35_rst = rst;
	assign branch_26_in2_data = fork_35__branch_26__data__0__anchor__in;
	assign fork_35__branch_26__data__0__anchor__out = fork_35_out1_data;
	assign branch_26_in2_valid = fork_35__branch_26__valid__0__anchor__in;
	assign fork_35__branch_26__valid__0__anchor__out = fork_35_out1_valid;
	assign fork_35_out1_ready = fork_35__branch_26__ready__0__anchor__in;
	assign fork_35__branch_26__ready__0__anchor__out = branch_26_in2_ready;
	assign branch_25_in2_data = fork_35__branch_25__data__0__anchor__in;
	assign fork_35__branch_25__data__0__anchor__out = fork_35_out2_data;
	assign branch_25_in2_valid = fork_35__branch_25__valid__0__anchor__in;
	assign fork_35__branch_25__valid__0__anchor__out = fork_35_out2_valid;
	assign fork_35_out2_ready = fork_35__branch_25__ready__0__anchor__in;
	assign fork_35__branch_25__ready__0__anchor__out = branch_25_in2_ready;
	assign branch_24_in2_data = fork_35__branch_24__data__0__anchor__in;
	assign fork_35__branch_24__data__0__anchor__out = fork_35_out3_data;
	assign branch_24_in2_valid = fork_35__branch_24__valid__0__anchor__in;
	assign fork_35__branch_24__valid__0__anchor__out = fork_35_out3_valid;
	assign fork_35_out3_ready = fork_35__branch_24__ready__0__anchor__in;
	assign fork_35__branch_24__ready__0__anchor__out = branch_24_in2_ready;
	assign branch_23_in2_data = fork_35__branch_23__data__0__anchor__in;
	assign fork_35__branch_23__data__0__anchor__out = fork_35_out4_data;
	assign branch_23_in2_valid = fork_35__branch_23__valid__0__anchor__in;
	assign fork_35__branch_23__valid__0__anchor__out = fork_35_out4_valid;
	assign fork_35_out4_ready = fork_35__branch_23__ready__0__anchor__in;
	assign fork_35__branch_23__ready__0__anchor__out = branch_23_in2_ready;
	assign branch_22_in2_data = fork_35__branch_22__data__0__anchor__in;
	assign fork_35__branch_22__data__0__anchor__out = fork_35_out5_data;
	assign branch_22_in2_valid = fork_35__branch_22__valid__0__anchor__in;
	assign fork_35__branch_22__valid__0__anchor__out = fork_35_out5_valid;
	assign fork_35_out5_ready = fork_35__branch_22__ready__0__anchor__in;
	assign fork_35__branch_22__ready__0__anchor__out = branch_22_in2_ready;
	assign branchC_52_in2_data = fork_35__branchC_52__data__0__anchor__in;
	assign fork_35__branchC_52__data__0__anchor__out = fork_35_out6_data;
	assign branchC_52_in2_valid = fork_35__branchC_52__valid__0__anchor__in;
	assign fork_35__branchC_52__valid__0__anchor__out = fork_35_out6_valid;
	assign fork_35_out6_ready = fork_35__branchC_52__ready__0__anchor__in;
	assign fork_35__branchC_52__ready__0__anchor__out = branchC_52_in2_ready;
	assign branch_27_clk = clk;
	assign branch_27_rst = rst;
	assign Buffer_13_in1_data = branch_27__Buffer_13__data__0__anchor__in;
	assign branch_27__Buffer_13__data__0__anchor__out = branch_27_out1_data;
	assign Buffer_13_in1_valid = branch_27__Buffer_13__valid__0__anchor__in;
	assign branch_27__Buffer_13__valid__0__anchor__out = branch_27_out1_valid;
	assign branch_27_out1_ready = branch_27__Buffer_13__ready__0__anchor__in;
	assign branch_27__Buffer_13__ready__0__anchor__out = Buffer_13_in1_ready;
	assign sink_18_in1_data = branch_27__sink_18__data__0__anchor__in;
	assign branch_27__sink_18__data__0__anchor__out = branch_27_out2_data;
	assign sink_18_in1_valid = branch_27__sink_18__valid__0__anchor__in;
	assign branch_27__sink_18__valid__0__anchor__out = branch_27_out2_valid;
	assign branch_27_out2_ready = branch_27__sink_18__ready__0__anchor__in;
	assign branch_27__sink_18__ready__0__anchor__out = sink_18_in1_ready;
	assign branch_28_clk = clk;
	assign branch_28_rst = rst;
	assign Buffer_9_in1_data = branch_28__Buffer_9__data__0__anchor__in;
	assign branch_28__Buffer_9__data__0__anchor__out = branch_28_out1_data;
	assign Buffer_9_in1_valid = branch_28__Buffer_9__valid__0__anchor__in;
	assign branch_28__Buffer_9__valid__0__anchor__out = branch_28_out1_valid;
	assign branch_28_out1_ready = branch_28__Buffer_9__ready__0__anchor__in;
	assign branch_28__Buffer_9__ready__0__anchor__out = Buffer_9_in1_ready;
	assign sink_19_in1_data = branch_28__sink_19__data__0__anchor__in;
	assign branch_28__sink_19__data__0__anchor__out = branch_28_out2_data;
	assign sink_19_in1_valid = branch_28__sink_19__valid__0__anchor__in;
	assign branch_28__sink_19__valid__0__anchor__out = branch_28_out2_valid;
	assign branch_28_out2_ready = branch_28__sink_19__ready__0__anchor__in;
	assign branch_28__sink_19__ready__0__anchor__out = sink_19_in1_ready;
	assign branch_29_clk = clk;
	assign branch_29_rst = rst;
	assign Buffer_24_in1_data = branch_29__Buffer_24__data__0__anchor__in;
	assign branch_29__Buffer_24__data__0__anchor__out = branch_29_out1_data;
	assign Buffer_24_in1_valid = branch_29__Buffer_24__valid__0__anchor__in;
	assign branch_29__Buffer_24__valid__0__anchor__out = branch_29_out1_valid;
	assign branch_29_out1_ready = branch_29__Buffer_24__ready__0__anchor__in;
	assign branch_29__Buffer_24__ready__0__anchor__out = Buffer_24_in1_ready;
	assign phi_n19_in1_data = branch_29__phi_n19__data__0__anchor__in;
	assign branch_29__phi_n19__data__0__anchor__out = branch_29_out2_data;
	assign phi_n19_in1_valid = branch_29__phi_n19__valid__0__anchor__in;
	assign branch_29__phi_n19__valid__0__anchor__out = branch_29_out2_valid;
	assign branch_29_out2_ready = branch_29__phi_n19__ready__0__anchor__in;
	assign branch_29__phi_n19__ready__0__anchor__out = phi_n19_in1_ready;
	assign fork_36_clk = clk;
	assign fork_36_rst = rst;
	assign branch_29_in2_data = fork_36__branch_29__data__0__anchor__in;
	assign fork_36__branch_29__data__0__anchor__out = fork_36_out1_data;
	assign branch_29_in2_valid = fork_36__branch_29__valid__0__anchor__in;
	assign fork_36__branch_29__valid__0__anchor__out = fork_36_out1_valid;
	assign fork_36_out1_ready = fork_36__branch_29__ready__0__anchor__in;
	assign fork_36__branch_29__ready__0__anchor__out = branch_29_in2_ready;
	assign branch_28_in2_data = fork_36__branch_28__data__0__anchor__in;
	assign fork_36__branch_28__data__0__anchor__out = fork_36_out2_data;
	assign branch_28_in2_valid = fork_36__branch_28__valid__0__anchor__in;
	assign fork_36__branch_28__valid__0__anchor__out = fork_36_out2_valid;
	assign fork_36_out2_ready = fork_36__branch_28__ready__0__anchor__in;
	assign fork_36__branch_28__ready__0__anchor__out = branch_28_in2_ready;
	assign branch_27_in2_data = fork_36__branch_27__data__0__anchor__in;
	assign fork_36__branch_27__data__0__anchor__out = fork_36_out3_data;
	assign branch_27_in2_valid = fork_36__branch_27__valid__0__anchor__in;
	assign fork_36__branch_27__valid__0__anchor__out = fork_36_out3_valid;
	assign fork_36_out3_ready = fork_36__branch_27__ready__0__anchor__in;
	assign fork_36__branch_27__ready__0__anchor__out = branch_27_in2_ready;
	assign branchC_53_in2_data = fork_36__branchC_53__data__0__anchor__in;
	assign fork_36__branchC_53__data__0__anchor__out = fork_36_out4_data;
	assign branchC_53_in2_valid = fork_36__branchC_53__valid__0__anchor__in;
	assign fork_36__branchC_53__valid__0__anchor__out = fork_36_out4_valid;
	assign fork_36_out4_ready = fork_36__branchC_53__ready__0__anchor__in;
	assign fork_36__branchC_53__ready__0__anchor__out = branchC_53_in2_ready;
	assign branch_30_clk = clk;
	assign branch_30_rst = rst;
	assign phi_63_in2_data = branch_30__phi_63__data__0__anchor__in;
	assign branch_30__phi_63__data__0__anchor__out = branch_30_out1_data;
	assign phi_63_in2_valid = branch_30__phi_63__valid__0__anchor__in;
	assign branch_30__phi_63__valid__0__anchor__out = branch_30_out1_valid;
	assign branch_30_out1_ready = branch_30__phi_63__ready__0__anchor__in;
	assign branch_30__phi_63__ready__0__anchor__out = phi_63_in2_ready;
	assign sink_20_in1_data = branch_30__sink_20__data__0__anchor__in;
	assign branch_30__sink_20__data__0__anchor__out = branch_30_out2_data;
	assign sink_20_in1_valid = branch_30__sink_20__valid__0__anchor__in;
	assign branch_30__sink_20__valid__0__anchor__out = branch_30_out2_valid;
	assign branch_30_out2_ready = branch_30__sink_20__ready__0__anchor__in;
	assign branch_30__sink_20__ready__0__anchor__out = sink_20_in1_ready;
	assign branch_31_clk = clk;
	assign branch_31_rst = rst;
	assign phi_n20_in1_data = branch_31__phi_n20__data__0__anchor__in;
	assign branch_31__phi_n20__data__0__anchor__out = branch_31_out1_data;
	assign phi_n20_in1_valid = branch_31__phi_n20__valid__0__anchor__in;
	assign branch_31__phi_n20__valid__0__anchor__out = branch_31_out1_valid;
	assign branch_31_out1_ready = branch_31__phi_n20__ready__0__anchor__in;
	assign branch_31__phi_n20__ready__0__anchor__out = phi_n20_in1_ready;
	assign sink_21_in1_data = branch_31__sink_21__data__0__anchor__in;
	assign branch_31__sink_21__data__0__anchor__out = branch_31_out2_data;
	assign sink_21_in1_valid = branch_31__sink_21__valid__0__anchor__in;
	assign branch_31__sink_21__valid__0__anchor__out = branch_31_out2_valid;
	assign branch_31_out2_ready = branch_31__sink_21__ready__0__anchor__in;
	assign branch_31__sink_21__ready__0__anchor__out = sink_21_in1_ready;
	assign fork_37_clk = clk;
	assign fork_37_rst = rst;
	assign branch_31_in2_data = fork_37__branch_31__data__0__anchor__in;
	assign fork_37__branch_31__data__0__anchor__out = fork_37_out1_data;
	assign branch_31_in2_valid = fork_37__branch_31__valid__0__anchor__in;
	assign fork_37__branch_31__valid__0__anchor__out = fork_37_out1_valid;
	assign fork_37_out1_ready = fork_37__branch_31__ready__0__anchor__in;
	assign fork_37__branch_31__ready__0__anchor__out = branch_31_in2_ready;
	assign branch_30_in2_data = fork_37__branch_30__data__0__anchor__in;
	assign fork_37__branch_30__data__0__anchor__out = fork_37_out2_data;
	assign branch_30_in2_valid = fork_37__branch_30__valid__0__anchor__in;
	assign fork_37__branch_30__valid__0__anchor__out = fork_37_out2_valid;
	assign fork_37_out2_ready = fork_37__branch_30__ready__0__anchor__in;
	assign fork_37__branch_30__ready__0__anchor__out = branch_30_in2_ready;
	assign branchC_54_in2_data = fork_37__branchC_54__data__0__anchor__in;
	assign fork_37__branchC_54__data__0__anchor__out = fork_37_out3_data;
	assign branchC_54_in2_valid = fork_37__branchC_54__valid__0__anchor__in;
	assign fork_37__branchC_54__valid__0__anchor__out = fork_37_out3_valid;
	assign fork_37_out3_ready = fork_37__branchC_54__ready__0__anchor__in;
	assign fork_37__branchC_54__ready__0__anchor__out = branchC_54_in2_ready;
	assign branch_32_clk = clk;
	assign branch_32_rst = rst;
	assign Buffer_10_in1_data = branch_32__Buffer_10__data__0__anchor__in;
	assign branch_32__Buffer_10__data__0__anchor__out = branch_32_out1_data;
	assign Buffer_10_in1_valid = branch_32__Buffer_10__valid__0__anchor__in;
	assign branch_32__Buffer_10__valid__0__anchor__out = branch_32_out1_valid;
	assign branch_32_out1_ready = branch_32__Buffer_10__ready__0__anchor__in;
	assign branch_32__Buffer_10__ready__0__anchor__out = Buffer_10_in1_ready;
	assign sink_22_in1_data = branch_32__sink_22__data__0__anchor__in;
	assign branch_32__sink_22__data__0__anchor__out = branch_32_out2_data;
	assign sink_22_in1_valid = branch_32__sink_22__valid__0__anchor__in;
	assign branch_32__sink_22__valid__0__anchor__out = branch_32_out2_valid;
	assign branch_32_out2_ready = branch_32__sink_22__ready__0__anchor__in;
	assign branch_32__sink_22__ready__0__anchor__out = sink_22_in1_ready;
	assign branch_33_clk = clk;
	assign branch_33_rst = rst;
	assign Buffer_28_in1_data = branch_33__Buffer_28__data__0__anchor__in;
	assign branch_33__Buffer_28__data__0__anchor__out = branch_33_out1_data;
	assign Buffer_28_in1_valid = branch_33__Buffer_28__valid__0__anchor__in;
	assign branch_33__Buffer_28__valid__0__anchor__out = branch_33_out1_valid;
	assign branch_33_out1_ready = branch_33__Buffer_28__ready__0__anchor__in;
	assign branch_33__Buffer_28__ready__0__anchor__out = Buffer_28_in1_ready;
	assign phi_n21_in1_data = branch_33__phi_n21__data__0__anchor__in;
	assign branch_33__phi_n21__data__0__anchor__out = branch_33_out2_data;
	assign phi_n21_in1_valid = branch_33__phi_n21__valid__0__anchor__in;
	assign branch_33__phi_n21__valid__0__anchor__out = branch_33_out2_valid;
	assign branch_33_out2_ready = branch_33__phi_n21__ready__0__anchor__in;
	assign branch_33__phi_n21__ready__0__anchor__out = phi_n21_in1_ready;
	assign fork_38_clk = clk;
	assign fork_38_rst = rst;
	assign branch_33_in2_data = fork_38__branch_33__data__0__anchor__in;
	assign fork_38__branch_33__data__0__anchor__out = fork_38_out1_data;
	assign branch_33_in2_valid = fork_38__branch_33__valid__0__anchor__in;
	assign fork_38__branch_33__valid__0__anchor__out = fork_38_out1_valid;
	assign fork_38_out1_ready = fork_38__branch_33__ready__0__anchor__in;
	assign fork_38__branch_33__ready__0__anchor__out = branch_33_in2_ready;
	assign branch_32_in2_data = fork_38__branch_32__data__0__anchor__in;
	assign fork_38__branch_32__data__0__anchor__out = fork_38_out2_data;
	assign branch_32_in2_valid = fork_38__branch_32__valid__0__anchor__in;
	assign fork_38__branch_32__valid__0__anchor__out = fork_38_out2_valid;
	assign fork_38_out2_ready = fork_38__branch_32__ready__0__anchor__in;
	assign fork_38__branch_32__ready__0__anchor__out = branch_32_in2_ready;
	assign branchC_55_in2_data = fork_38__branchC_55__data__0__anchor__in;
	assign fork_38__branchC_55__data__0__anchor__out = fork_38_out3_data;
	assign branchC_55_in2_valid = fork_38__branchC_55__valid__0__anchor__in;
	assign fork_38__branchC_55__valid__0__anchor__out = fork_38_out3_valid;
	assign fork_38_out3_ready = fork_38__branchC_55__ready__0__anchor__in;
	assign fork_38__branchC_55__ready__0__anchor__out = branchC_55_in2_ready;
	assign branch_34_clk = clk;
	assign branch_34_rst = rst;
	assign phi_77_in2_data = branch_34__phi_77__data__0__anchor__in;
	assign branch_34__phi_77__data__0__anchor__out = branch_34_out1_data;
	assign phi_77_in2_valid = branch_34__phi_77__valid__0__anchor__in;
	assign branch_34__phi_77__valid__0__anchor__out = branch_34_out1_valid;
	assign branch_34_out1_ready = branch_34__phi_77__ready__0__anchor__in;
	assign branch_34__phi_77__ready__0__anchor__out = phi_77_in2_ready;
	assign sink_23_in1_data = branch_34__sink_23__data__0__anchor__in;
	assign branch_34__sink_23__data__0__anchor__out = branch_34_out2_data;
	assign sink_23_in1_valid = branch_34__sink_23__valid__0__anchor__in;
	assign branch_34__sink_23__valid__0__anchor__out = branch_34_out2_valid;
	assign branch_34_out2_ready = branch_34__sink_23__ready__0__anchor__in;
	assign branch_34__sink_23__ready__0__anchor__out = sink_23_in1_ready;
	assign branch_35_clk = clk;
	assign branch_35_rst = rst;
	assign phi_n22_in1_data = branch_35__phi_n22__data__0__anchor__in;
	assign branch_35__phi_n22__data__0__anchor__out = branch_35_out1_data;
	assign phi_n22_in1_valid = branch_35__phi_n22__valid__0__anchor__in;
	assign branch_35__phi_n22__valid__0__anchor__out = branch_35_out1_valid;
	assign branch_35_out1_ready = branch_35__phi_n22__ready__0__anchor__in;
	assign branch_35__phi_n22__ready__0__anchor__out = phi_n22_in1_ready;
	assign sink_24_in1_data = branch_35__sink_24__data__0__anchor__in;
	assign branch_35__sink_24__data__0__anchor__out = branch_35_out2_data;
	assign sink_24_in1_valid = branch_35__sink_24__valid__0__anchor__in;
	assign branch_35__sink_24__valid__0__anchor__out = branch_35_out2_valid;
	assign branch_35_out2_ready = branch_35__sink_24__ready__0__anchor__in;
	assign branch_35__sink_24__ready__0__anchor__out = sink_24_in1_ready;
	assign fork_39_clk = clk;
	assign fork_39_rst = rst;
	assign branch_35_in2_data = fork_39__branch_35__data__0__anchor__in;
	assign fork_39__branch_35__data__0__anchor__out = fork_39_out1_data;
	assign branch_35_in2_valid = fork_39__branch_35__valid__0__anchor__in;
	assign fork_39__branch_35__valid__0__anchor__out = fork_39_out1_valid;
	assign fork_39_out1_ready = fork_39__branch_35__ready__0__anchor__in;
	assign fork_39__branch_35__ready__0__anchor__out = branch_35_in2_ready;
	assign branch_34_in2_data = fork_39__branch_34__data__0__anchor__in;
	assign fork_39__branch_34__data__0__anchor__out = fork_39_out2_data;
	assign branch_34_in2_valid = fork_39__branch_34__valid__0__anchor__in;
	assign fork_39__branch_34__valid__0__anchor__out = fork_39_out2_valid;
	assign fork_39_out2_ready = fork_39__branch_34__ready__0__anchor__in;
	assign fork_39__branch_34__ready__0__anchor__out = branch_34_in2_ready;
	assign branchC_56_in2_data = fork_39__branchC_56__data__0__anchor__in;
	assign fork_39__branchC_56__data__0__anchor__out = fork_39_out3_data;
	assign branchC_56_in2_valid = fork_39__branchC_56__valid__0__anchor__in;
	assign fork_39__branchC_56__valid__0__anchor__out = fork_39_out3_valid;
	assign fork_39_out3_ready = fork_39__branchC_56__ready__0__anchor__in;
	assign fork_39__branchC_56__ready__0__anchor__out = branchC_56_in2_ready;
	assign branch_36_clk = clk;
	assign branch_36_rst = rst;
	assign phi_82_in2_data = branch_36__phi_82__data__0__anchor__in;
	assign branch_36__phi_82__data__0__anchor__out = branch_36_out1_data;
	assign phi_82_in2_valid = branch_36__phi_82__valid__0__anchor__in;
	assign branch_36__phi_82__valid__0__anchor__out = branch_36_out1_valid;
	assign branch_36_out1_ready = branch_36__phi_82__ready__0__anchor__in;
	assign branch_36__phi_82__ready__0__anchor__out = phi_82_in2_ready;
	assign sink_25_in1_data = branch_36__sink_25__data__0__anchor__in;
	assign branch_36__sink_25__data__0__anchor__out = branch_36_out2_data;
	assign sink_25_in1_valid = branch_36__sink_25__valid__0__anchor__in;
	assign branch_36__sink_25__valid__0__anchor__out = branch_36_out2_valid;
	assign branch_36_out2_ready = branch_36__sink_25__ready__0__anchor__in;
	assign branch_36__sink_25__ready__0__anchor__out = sink_25_in1_ready;
	assign branch_37_clk = clk;
	assign branch_37_rst = rst;
	assign phi_83_in2_data = branch_37__phi_83__data__0__anchor__in;
	assign branch_37__phi_83__data__0__anchor__out = branch_37_out1_data;
	assign phi_83_in2_valid = branch_37__phi_83__valid__0__anchor__in;
	assign branch_37__phi_83__valid__0__anchor__out = branch_37_out1_valid;
	assign branch_37_out1_ready = branch_37__phi_83__ready__0__anchor__in;
	assign branch_37__phi_83__ready__0__anchor__out = phi_83_in2_ready;
	assign sink_26_in1_data = branch_37__sink_26__data__0__anchor__in;
	assign branch_37__sink_26__data__0__anchor__out = branch_37_out2_data;
	assign sink_26_in1_valid = branch_37__sink_26__valid__0__anchor__in;
	assign branch_37__sink_26__valid__0__anchor__out = branch_37_out2_valid;
	assign branch_37_out2_ready = branch_37__sink_26__ready__0__anchor__in;
	assign branch_37__sink_26__ready__0__anchor__out = sink_26_in1_ready;
	assign branch_38_clk = clk;
	assign branch_38_rst = rst;
	assign phi_n27_in1_data = branch_38__phi_n27__data__0__anchor__in;
	assign branch_38__phi_n27__data__0__anchor__out = branch_38_out1_data;
	assign phi_n27_in1_valid = branch_38__phi_n27__valid__0__anchor__in;
	assign branch_38__phi_n27__valid__0__anchor__out = branch_38_out1_valid;
	assign branch_38_out1_ready = branch_38__phi_n27__ready__0__anchor__in;
	assign branch_38__phi_n27__ready__0__anchor__out = phi_n27_in1_ready;
	assign sink_27_in1_data = branch_38__sink_27__data__0__anchor__in;
	assign branch_38__sink_27__data__0__anchor__out = branch_38_out2_data;
	assign sink_27_in1_valid = branch_38__sink_27__valid__0__anchor__in;
	assign branch_38__sink_27__valid__0__anchor__out = branch_38_out2_valid;
	assign branch_38_out2_ready = branch_38__sink_27__ready__0__anchor__in;
	assign branch_38__sink_27__ready__0__anchor__out = sink_27_in1_ready;
	assign branch_39_clk = clk;
	assign branch_39_rst = rst;
	assign phi_n26_in1_data = branch_39__phi_n26__data__0__anchor__in;
	assign branch_39__phi_n26__data__0__anchor__out = branch_39_out1_data;
	assign phi_n26_in1_valid = branch_39__phi_n26__valid__0__anchor__in;
	assign branch_39__phi_n26__valid__0__anchor__out = branch_39_out1_valid;
	assign branch_39_out1_ready = branch_39__phi_n26__ready__0__anchor__in;
	assign branch_39__phi_n26__ready__0__anchor__out = phi_n26_in1_ready;
	assign sink_28_in1_data = branch_39__sink_28__data__0__anchor__in;
	assign branch_39__sink_28__data__0__anchor__out = branch_39_out2_data;
	assign sink_28_in1_valid = branch_39__sink_28__valid__0__anchor__in;
	assign branch_39__sink_28__valid__0__anchor__out = branch_39_out2_valid;
	assign branch_39_out2_ready = branch_39__sink_28__ready__0__anchor__in;
	assign branch_39__sink_28__ready__0__anchor__out = sink_28_in1_ready;
	assign fork_40_clk = clk;
	assign fork_40_rst = rst;
	assign branch_39_in2_data = fork_40__branch_39__data__0__anchor__in;
	assign fork_40__branch_39__data__0__anchor__out = fork_40_out1_data;
	assign branch_39_in2_valid = fork_40__branch_39__valid__0__anchor__in;
	assign fork_40__branch_39__valid__0__anchor__out = fork_40_out1_valid;
	assign fork_40_out1_ready = fork_40__branch_39__ready__0__anchor__in;
	assign fork_40__branch_39__ready__0__anchor__out = branch_39_in2_ready;
	assign branch_38_in2_data = fork_40__branch_38__data__0__anchor__in;
	assign fork_40__branch_38__data__0__anchor__out = fork_40_out2_data;
	assign branch_38_in2_valid = fork_40__branch_38__valid__0__anchor__in;
	assign fork_40__branch_38__valid__0__anchor__out = fork_40_out2_valid;
	assign fork_40_out2_ready = fork_40__branch_38__ready__0__anchor__in;
	assign fork_40__branch_38__ready__0__anchor__out = branch_38_in2_ready;
	assign branch_37_in2_data = fork_40__branch_37__data__0__anchor__in;
	assign fork_40__branch_37__data__0__anchor__out = fork_40_out3_data;
	assign branch_37_in2_valid = fork_40__branch_37__valid__0__anchor__in;
	assign fork_40__branch_37__valid__0__anchor__out = fork_40_out3_valid;
	assign fork_40_out3_ready = fork_40__branch_37__ready__0__anchor__in;
	assign fork_40__branch_37__ready__0__anchor__out = branch_37_in2_ready;
	assign branch_36_in2_data = fork_40__branch_36__data__0__anchor__in;
	assign fork_40__branch_36__data__0__anchor__out = fork_40_out4_data;
	assign branch_36_in2_valid = fork_40__branch_36__valid__0__anchor__in;
	assign fork_40__branch_36__valid__0__anchor__out = fork_40_out4_valid;
	assign fork_40_out4_ready = fork_40__branch_36__ready__0__anchor__in;
	assign fork_40__branch_36__ready__0__anchor__out = branch_36_in2_ready;
	assign branchC_57_in2_data = fork_40__branchC_57__data__0__anchor__in;
	assign fork_40__branchC_57__data__0__anchor__out = fork_40_out5_data;
	assign branchC_57_in2_valid = fork_40__branchC_57__valid__0__anchor__in;
	assign fork_40__branchC_57__valid__0__anchor__out = fork_40_out5_valid;
	assign fork_40_out5_ready = fork_40__branchC_57__ready__0__anchor__in;
	assign fork_40__branchC_57__ready__0__anchor__out = branchC_57_in2_ready;
	assign branch_40_clk = clk;
	assign branch_40_rst = rst;
	assign Buffer_8_in1_data = branch_40__Buffer_8__data__0__anchor__in;
	assign branch_40__Buffer_8__data__0__anchor__out = branch_40_out1_data;
	assign Buffer_8_in1_valid = branch_40__Buffer_8__valid__0__anchor__in;
	assign branch_40__Buffer_8__valid__0__anchor__out = branch_40_out1_valid;
	assign branch_40_out1_ready = branch_40__Buffer_8__ready__0__anchor__in;
	assign branch_40__Buffer_8__ready__0__anchor__out = Buffer_8_in1_ready;
	assign phi_n23_in1_data = branch_40__phi_n23__data__0__anchor__in;
	assign branch_40__phi_n23__data__0__anchor__out = branch_40_out2_data;
	assign phi_n23_in1_valid = branch_40__phi_n23__valid__0__anchor__in;
	assign branch_40__phi_n23__valid__0__anchor__out = branch_40_out2_valid;
	assign branch_40_out2_ready = branch_40__phi_n23__ready__0__anchor__in;
	assign branch_40__phi_n23__ready__0__anchor__out = phi_n23_in1_ready;
	assign branch_41_clk = clk;
	assign branch_41_rst = rst;
	assign Buffer_29_in1_data = branch_41__Buffer_29__data__0__anchor__in;
	assign branch_41__Buffer_29__data__0__anchor__out = branch_41_out1_data;
	assign Buffer_29_in1_valid = branch_41__Buffer_29__valid__0__anchor__in;
	assign branch_41__Buffer_29__valid__0__anchor__out = branch_41_out1_valid;
	assign branch_41_out1_ready = branch_41__Buffer_29__ready__0__anchor__in;
	assign branch_41__Buffer_29__ready__0__anchor__out = Buffer_29_in1_ready;
	assign sink_29_in1_data = branch_41__sink_29__data__0__anchor__in;
	assign branch_41__sink_29__data__0__anchor__out = branch_41_out2_data;
	assign sink_29_in1_valid = branch_41__sink_29__valid__0__anchor__in;
	assign branch_41__sink_29__valid__0__anchor__out = branch_41_out2_valid;
	assign branch_41_out2_ready = branch_41__sink_29__ready__0__anchor__in;
	assign branch_41__sink_29__ready__0__anchor__out = sink_29_in1_ready;
	assign branch_42_clk = clk;
	assign branch_42_rst = rst;
	assign Buffer_15_in1_data = branch_42__Buffer_15__data__0__anchor__in;
	assign branch_42__Buffer_15__data__0__anchor__out = branch_42_out1_data;
	assign Buffer_15_in1_valid = branch_42__Buffer_15__valid__0__anchor__in;
	assign branch_42__Buffer_15__valid__0__anchor__out = branch_42_out1_valid;
	assign branch_42_out1_ready = branch_42__Buffer_15__ready__0__anchor__in;
	assign branch_42__Buffer_15__ready__0__anchor__out = Buffer_15_in1_ready;
	assign phi_n24_in1_data = branch_42__phi_n24__data__0__anchor__in;
	assign branch_42__phi_n24__data__0__anchor__out = branch_42_out2_data;
	assign phi_n24_in1_valid = branch_42__phi_n24__valid__0__anchor__in;
	assign branch_42__phi_n24__valid__0__anchor__out = branch_42_out2_valid;
	assign branch_42_out2_ready = branch_42__phi_n24__ready__0__anchor__in;
	assign branch_42__phi_n24__ready__0__anchor__out = phi_n24_in1_ready;
	assign branch_43_clk = clk;
	assign branch_43_rst = rst;
	assign Buffer_23_in1_data = branch_43__Buffer_23__data__0__anchor__in;
	assign branch_43__Buffer_23__data__0__anchor__out = branch_43_out1_data;
	assign Buffer_23_in1_valid = branch_43__Buffer_23__valid__0__anchor__in;
	assign branch_43__Buffer_23__valid__0__anchor__out = branch_43_out1_valid;
	assign branch_43_out1_ready = branch_43__Buffer_23__ready__0__anchor__in;
	assign branch_43__Buffer_23__ready__0__anchor__out = Buffer_23_in1_ready;
	assign phi_n25_in1_data = branch_43__phi_n25__data__0__anchor__in;
	assign branch_43__phi_n25__data__0__anchor__out = branch_43_out2_data;
	assign phi_n25_in1_valid = branch_43__phi_n25__valid__0__anchor__in;
	assign branch_43__phi_n25__valid__0__anchor__out = branch_43_out2_valid;
	assign branch_43_out2_ready = branch_43__phi_n25__ready__0__anchor__in;
	assign branch_43__phi_n25__ready__0__anchor__out = phi_n25_in1_ready;
	assign fork_41_clk = clk;
	assign fork_41_rst = rst;
	assign branch_43_in2_data = fork_41__branch_43__data__0__anchor__in;
	assign fork_41__branch_43__data__0__anchor__out = fork_41_out1_data;
	assign branch_43_in2_valid = fork_41__branch_43__valid__0__anchor__in;
	assign fork_41__branch_43__valid__0__anchor__out = fork_41_out1_valid;
	assign fork_41_out1_ready = fork_41__branch_43__ready__0__anchor__in;
	assign fork_41__branch_43__ready__0__anchor__out = branch_43_in2_ready;
	assign branch_42_in2_data = fork_41__branch_42__data__0__anchor__in;
	assign fork_41__branch_42__data__0__anchor__out = fork_41_out2_data;
	assign branch_42_in2_valid = fork_41__branch_42__valid__0__anchor__in;
	assign fork_41__branch_42__valid__0__anchor__out = fork_41_out2_valid;
	assign fork_41_out2_ready = fork_41__branch_42__ready__0__anchor__in;
	assign fork_41__branch_42__ready__0__anchor__out = branch_42_in2_ready;
	assign branch_41_in2_data = fork_41__branch_41__data__0__anchor__in;
	assign fork_41__branch_41__data__0__anchor__out = fork_41_out3_data;
	assign branch_41_in2_valid = fork_41__branch_41__valid__0__anchor__in;
	assign fork_41__branch_41__valid__0__anchor__out = fork_41_out3_valid;
	assign fork_41_out3_ready = fork_41__branch_41__ready__0__anchor__in;
	assign fork_41__branch_41__ready__0__anchor__out = branch_41_in2_ready;
	assign branch_40_in2_data = fork_41__branch_40__data__0__anchor__in;
	assign fork_41__branch_40__data__0__anchor__out = fork_41_out4_data;
	assign branch_40_in2_valid = fork_41__branch_40__valid__0__anchor__in;
	assign fork_41__branch_40__valid__0__anchor__out = fork_41_out4_valid;
	assign fork_41_out4_ready = fork_41__branch_40__ready__0__anchor__in;
	assign fork_41__branch_40__ready__0__anchor__out = branch_40_in2_ready;
	assign branchC_58_in2_data = fork_41__branchC_58__data__0__anchor__in;
	assign fork_41__branchC_58__data__0__anchor__out = fork_41_out5_data;
	assign branchC_58_in2_valid = fork_41__branchC_58__valid__0__anchor__in;
	assign fork_41__branchC_58__valid__0__anchor__out = fork_41_out5_valid;
	assign fork_41_out5_ready = fork_41__branchC_58__ready__0__anchor__in;
	assign fork_41__branchC_58__ready__0__anchor__out = branchC_58_in2_ready;
	assign branch_44_clk = clk;
	assign branch_44_rst = rst;
	assign Buffer_11_in1_data = branch_44__Buffer_11__data__0__anchor__in;
	assign branch_44__Buffer_11__data__0__anchor__out = branch_44_out1_data;
	assign Buffer_11_in1_valid = branch_44__Buffer_11__valid__0__anchor__in;
	assign branch_44__Buffer_11__valid__0__anchor__out = branch_44_out1_valid;
	assign branch_44_out1_ready = branch_44__Buffer_11__ready__0__anchor__in;
	assign branch_44__Buffer_11__ready__0__anchor__out = Buffer_11_in1_ready;
	assign sink_30_in1_data = branch_44__sink_30__data__0__anchor__in;
	assign branch_44__sink_30__data__0__anchor__out = branch_44_out2_data;
	assign sink_30_in1_valid = branch_44__sink_30__valid__0__anchor__in;
	assign branch_44__sink_30__valid__0__anchor__out = branch_44_out2_valid;
	assign branch_44_out2_ready = branch_44__sink_30__ready__0__anchor__in;
	assign branch_44__sink_30__ready__0__anchor__out = sink_30_in1_ready;
	assign branch_45_clk = clk;
	assign branch_45_rst = rst;
	assign Buffer_0_in1_data = branch_45__Buffer_0__data__0__anchor__in;
	assign branch_45__Buffer_0__data__0__anchor__out = branch_45_out1_data;
	assign Buffer_0_in1_valid = branch_45__Buffer_0__valid__0__anchor__in;
	assign branch_45__Buffer_0__valid__0__anchor__out = branch_45_out1_valid;
	assign branch_45_out1_ready = branch_45__Buffer_0__ready__0__anchor__in;
	assign branch_45__Buffer_0__ready__0__anchor__out = Buffer_0_in1_ready;
	assign sink_31_in1_data = branch_45__sink_31__data__0__anchor__in;
	assign branch_45__sink_31__data__0__anchor__out = branch_45_out2_data;
	assign sink_31_in1_valid = branch_45__sink_31__valid__0__anchor__in;
	assign branch_45__sink_31__valid__0__anchor__out = branch_45_out2_valid;
	assign branch_45_out2_ready = branch_45__sink_31__ready__0__anchor__in;
	assign branch_45__sink_31__ready__0__anchor__out = sink_31_in1_ready;
	assign fork_42_clk = clk;
	assign fork_42_rst = rst;
	assign branch_45_in2_data = fork_42__branch_45__data__0__anchor__in;
	assign fork_42__branch_45__data__0__anchor__out = fork_42_out1_data;
	assign branch_45_in2_valid = fork_42__branch_45__valid__0__anchor__in;
	assign fork_42__branch_45__valid__0__anchor__out = fork_42_out1_valid;
	assign fork_42_out1_ready = fork_42__branch_45__ready__0__anchor__in;
	assign fork_42__branch_45__ready__0__anchor__out = branch_45_in2_ready;
	assign branch_44_in2_data = fork_42__branch_44__data__0__anchor__in;
	assign fork_42__branch_44__data__0__anchor__out = fork_42_out2_data;
	assign branch_44_in2_valid = fork_42__branch_44__valid__0__anchor__in;
	assign fork_42__branch_44__valid__0__anchor__out = fork_42_out2_valid;
	assign fork_42_out2_ready = fork_42__branch_44__ready__0__anchor__in;
	assign fork_42__branch_44__ready__0__anchor__out = branch_44_in2_ready;
	assign branchC_59_in2_data = fork_42__branchC_59__data__0__anchor__in;
	assign fork_42__branchC_59__data__0__anchor__out = fork_42_out3_data;
	assign branchC_59_in2_valid = fork_42__branchC_59__valid__0__anchor__in;
	assign fork_42__branchC_59__valid__0__anchor__out = fork_42_out3_valid;
	assign fork_42_out3_ready = fork_42__branchC_59__ready__0__anchor__in;
	assign fork_42__branchC_59__ready__0__anchor__out = branchC_59_in2_ready;
	assign MC_A_clk = clk;
	assign MC_A_rst = rst;
	assign A_ce0 = A_we0;
	assign load_8_in1_data = MC_A__load_8__data__0__anchor__in;
	assign MC_A__load_8__data__0__anchor__out = MC_A_out1_data;
	assign load_8_in1_valid = MC_A__load_8__valid__0__anchor__in;
	assign MC_A__load_8__valid__0__anchor__out = MC_A_out1_valid;
	assign MC_A_out1_ready = MC_A__load_8__ready__0__anchor__in;
	assign MC_A__load_8__ready__0__anchor__out = load_8_in1_ready;
	assign load_47_in1_data = MC_A__load_47__data__0__anchor__in;
	assign MC_A__load_47__data__0__anchor__out = MC_A_out2_data;
	assign load_47_in1_valid = MC_A__load_47__valid__0__anchor__in;
	assign MC_A__load_47__valid__0__anchor__out = MC_A_out2_valid;
	assign MC_A_out2_ready = MC_A__load_47__ready__0__anchor__in;
	assign MC_A__load_47__ready__0__anchor__out = load_47_in1_ready;
	assign load_88_in1_data = MC_A__load_88__data__0__anchor__in;
	assign MC_A__load_88__data__0__anchor__out = MC_A_out3_data;
	assign load_88_in1_valid = MC_A__load_88__valid__0__anchor__in;
	assign MC_A__load_88__valid__0__anchor__out = MC_A_out3_valid;
	assign MC_A_out3_ready = MC_A__load_88__ready__0__anchor__in;
	assign MC_A__load_88__ready__0__anchor__out = load_88_in1_ready;
	assign end_0_in1_data = MC_A__end_0__data__0__anchor__in;
	assign MC_A__end_0__data__0__anchor__out = MC_A_out4_data;
	assign end_0_in1_valid = MC_A__end_0__valid__0__anchor__in;
	assign MC_A__end_0__valid__0__anchor__out = MC_A_out4_valid;
	assign MC_A_out4_ready = MC_A__end_0__ready__0__anchor__in;
	assign MC_A__end_0__ready__0__anchor__out = end_0_in1_ready;
	assign MC_u1_clk = clk;
	assign MC_u1_rst = rst;
	assign u1_ce0 = u1_we0;
	assign MC_u1_in2_valid = 0;
	assign MC_u1_in2_data = 0;
	assign load_11_in1_data = MC_u1__load_11__data__0__anchor__in;
	assign MC_u1__load_11__data__0__anchor__out = MC_u1_out1_data;
	assign load_11_in1_valid = MC_u1__load_11__valid__0__anchor__in;
	assign MC_u1__load_11__valid__0__anchor__out = MC_u1_out1_valid;
	assign MC_u1_out1_ready = MC_u1__load_11__ready__0__anchor__in;
	assign MC_u1__load_11__ready__0__anchor__out = load_11_in1_ready;
	assign end_0_in2_data = MC_u1__end_0__data__0__anchor__in;
	assign MC_u1__end_0__data__0__anchor__out = MC_u1_out2_data;
	assign end_0_in2_valid = MC_u1__end_0__valid__0__anchor__in;
	assign MC_u1__end_0__valid__0__anchor__out = MC_u1_out2_valid;
	assign MC_u1_out2_ready = MC_u1__end_0__ready__0__anchor__in;
	assign MC_u1__end_0__ready__0__anchor__out = end_0_in2_ready;
	assign MC_v1_clk = clk;
	assign MC_v1_rst = rst;
	assign v1_ce0 = v1_we0;
	assign MC_v1_in2_valid = 0;
	assign MC_v1_in2_data = 0;
	assign load_14_in1_data = MC_v1__load_14__data__0__anchor__in;
	assign MC_v1__load_14__data__0__anchor__out = MC_v1_out1_data;
	assign load_14_in1_valid = MC_v1__load_14__valid__0__anchor__in;
	assign MC_v1__load_14__valid__0__anchor__out = MC_v1_out1_valid;
	assign MC_v1_out1_ready = MC_v1__load_14__ready__0__anchor__in;
	assign MC_v1__load_14__ready__0__anchor__out = load_14_in1_ready;
	assign end_0_in3_data = MC_v1__end_0__data__0__anchor__in;
	assign MC_v1__end_0__data__0__anchor__out = MC_v1_out2_data;
	assign end_0_in3_valid = MC_v1__end_0__valid__0__anchor__in;
	assign MC_v1__end_0__valid__0__anchor__out = MC_v1_out2_valid;
	assign MC_v1_out2_ready = MC_v1__end_0__ready__0__anchor__in;
	assign MC_v1__end_0__ready__0__anchor__out = end_0_in3_ready;
	assign MC_u2_clk = clk;
	assign MC_u2_rst = rst;
	assign u2_ce0 = u2_we0;
	assign MC_u2_in2_valid = 0;
	assign MC_u2_in2_data = 0;
	assign load_19_in1_data = MC_u2__load_19__data__0__anchor__in;
	assign MC_u2__load_19__data__0__anchor__out = MC_u2_out1_data;
	assign load_19_in1_valid = MC_u2__load_19__valid__0__anchor__in;
	assign MC_u2__load_19__valid__0__anchor__out = MC_u2_out1_valid;
	assign MC_u2_out1_ready = MC_u2__load_19__ready__0__anchor__in;
	assign MC_u2__load_19__ready__0__anchor__out = load_19_in1_ready;
	assign end_0_in4_data = MC_u2__end_0__data__0__anchor__in;
	assign MC_u2__end_0__data__0__anchor__out = MC_u2_out2_data;
	assign end_0_in4_valid = MC_u2__end_0__valid__0__anchor__in;
	assign MC_u2__end_0__valid__0__anchor__out = MC_u2_out2_valid;
	assign MC_u2_out2_ready = MC_u2__end_0__ready__0__anchor__in;
	assign MC_u2__end_0__ready__0__anchor__out = end_0_in4_ready;
	assign MC_v2_clk = clk;
	assign MC_v2_rst = rst;
	assign v2_ce0 = v2_we0;
	assign MC_v2_in2_valid = 0;
	assign MC_v2_in2_data = 0;
	assign load_22_in1_data = MC_v2__load_22__data__0__anchor__in;
	assign MC_v2__load_22__data__0__anchor__out = MC_v2_out1_data;
	assign load_22_in1_valid = MC_v2__load_22__valid__0__anchor__in;
	assign MC_v2__load_22__valid__0__anchor__out = MC_v2_out1_valid;
	assign MC_v2_out1_ready = MC_v2__load_22__ready__0__anchor__in;
	assign MC_v2__load_22__ready__0__anchor__out = load_22_in1_ready;
	assign end_0_in5_data = MC_v2__end_0__data__0__anchor__in;
	assign MC_v2__end_0__data__0__anchor__out = MC_v2_out2_data;
	assign end_0_in5_valid = MC_v2__end_0__valid__0__anchor__in;
	assign MC_v2__end_0__valid__0__anchor__out = MC_v2_out2_valid;
	assign MC_v2_out2_ready = MC_v2__end_0__ready__0__anchor__in;
	assign MC_v2__end_0__ready__0__anchor__out = end_0_in5_ready;
	assign cst_25_clk = clk;
	assign cst_25_rst = rst;
	assign MC_A_in1_data = cst_25__MC_A__data__0__anchor__in;
	assign cst_25__MC_A__data__0__anchor__out = cst_25_out1_data;
	assign MC_A_in1_valid = cst_25__MC_A__valid__0__anchor__in;
	assign cst_25__MC_A__valid__0__anchor__out = cst_25_out1_valid;
	assign cst_25_out1_ready = cst_25__MC_A__ready__0__anchor__in;
	assign cst_25__MC_A__ready__0__anchor__out = MC_A_in1_ready;
	assign MC_x_clk = clk;
	assign MC_x_rst = rst;
	assign x_ce0 = x_we0;
	assign load_39_in1_data = MC_x__load_39__data__0__anchor__in;
	assign MC_x__load_39__data__0__anchor__out = MC_x_out1_data;
	assign load_39_in1_valid = MC_x__load_39__valid__0__anchor__in;
	assign MC_x__load_39__valid__0__anchor__out = MC_x_out1_valid;
	assign MC_x_out1_ready = MC_x__load_39__ready__0__anchor__in;
	assign MC_x__load_39__ready__0__anchor__out = load_39_in1_ready;
	assign load_66_in1_data = MC_x__load_66__data__0__anchor__in;
	assign MC_x__load_66__data__0__anchor__out = MC_x_out2_data;
	assign load_66_in1_valid = MC_x__load_66__valid__0__anchor__in;
	assign MC_x__load_66__valid__0__anchor__out = MC_x_out2_valid;
	assign MC_x_out2_ready = MC_x__load_66__ready__0__anchor__in;
	assign MC_x__load_66__ready__0__anchor__out = load_66_in1_ready;
	assign load_92_in1_data = MC_x__load_92__data__0__anchor__in;
	assign MC_x__load_92__data__0__anchor__out = MC_x_out3_data;
	assign load_92_in1_valid = MC_x__load_92__valid__0__anchor__in;
	assign MC_x__load_92__valid__0__anchor__out = MC_x_out3_valid;
	assign MC_x_out3_ready = MC_x__load_92__ready__0__anchor__in;
	assign MC_x__load_92__ready__0__anchor__out = load_92_in1_ready;
	assign end_0_in6_data = MC_x__end_0__data__0__anchor__in;
	assign MC_x__end_0__data__0__anchor__out = MC_x_out4_data;
	assign end_0_in6_valid = MC_x__end_0__valid__0__anchor__in;
	assign MC_x__end_0__valid__0__anchor__out = MC_x_out4_valid;
	assign MC_x_out4_ready = MC_x__end_0__ready__0__anchor__in;
	assign MC_x__end_0__ready__0__anchor__out = end_0_in6_ready;
	assign MC_y_clk = clk;
	assign MC_y_rst = rst;
	assign y_ce0 = y_we0;
	assign MC_y_in2_valid = 0;
	assign MC_y_in2_data = 0;
	assign load_51_in1_data = MC_y__load_51__data__0__anchor__in;
	assign MC_y__load_51__data__0__anchor__out = MC_y_out1_data;
	assign load_51_in1_valid = MC_y__load_51__valid__0__anchor__in;
	assign MC_y__load_51__valid__0__anchor__out = MC_y_out1_valid;
	assign MC_y_out1_ready = MC_y__load_51__ready__0__anchor__in;
	assign MC_y__load_51__ready__0__anchor__out = load_51_in1_ready;
	assign end_0_in7_data = MC_y__end_0__data__0__anchor__in;
	assign MC_y__end_0__data__0__anchor__out = MC_y_out2_data;
	assign end_0_in7_valid = MC_y__end_0__valid__0__anchor__in;
	assign MC_y__end_0__valid__0__anchor__out = MC_y_out2_valid;
	assign MC_y_out2_ready = MC_y__end_0__ready__0__anchor__in;
	assign MC_y__end_0__ready__0__anchor__out = end_0_in7_ready;
	assign cst_26_clk = clk;
	assign cst_26_rst = rst;
	assign MC_x_in1_data = cst_26__MC_x__data__0__anchor__in;
	assign cst_26__MC_x__data__0__anchor__out = cst_26_out1_data;
	assign MC_x_in1_valid = cst_26__MC_x__valid__0__anchor__in;
	assign cst_26__MC_x__valid__0__anchor__out = cst_26_out1_valid;
	assign cst_26_out1_ready = cst_26__MC_x__ready__0__anchor__in;
	assign cst_26__MC_x__ready__0__anchor__out = MC_x_in1_ready;
	assign MC_z_clk = clk;
	assign MC_z_rst = rst;
	assign z_ce0 = z_we0;
	assign MC_z_in2_valid = 0;
	assign MC_z_in2_data = 0;
	assign load_69_in1_data = MC_z__load_69__data__0__anchor__in;
	assign MC_z__load_69__data__0__anchor__out = MC_z_out1_data;
	assign load_69_in1_valid = MC_z__load_69__valid__0__anchor__in;
	assign MC_z__load_69__valid__0__anchor__out = MC_z_out1_valid;
	assign MC_z_out1_ready = MC_z__load_69__ready__0__anchor__in;
	assign MC_z__load_69__ready__0__anchor__out = load_69_in1_ready;
	assign end_0_in8_data = MC_z__end_0__data__0__anchor__in;
	assign MC_z__end_0__data__0__anchor__out = MC_z_out2_data;
	assign end_0_in8_valid = MC_z__end_0__valid__0__anchor__in;
	assign MC_z__end_0__valid__0__anchor__out = MC_z_out2_valid;
	assign MC_z_out2_ready = MC_z__end_0__ready__0__anchor__in;
	assign MC_z__end_0__ready__0__anchor__out = end_0_in8_ready;
	assign cst_27_clk = clk;
	assign cst_27_rst = rst;
	assign MC_x_in2_data = cst_27__MC_x__data__0__anchor__in;
	assign cst_27__MC_x__data__0__anchor__out = cst_27_out1_data;
	assign MC_x_in2_valid = cst_27__MC_x__valid__0__anchor__in;
	assign cst_27__MC_x__valid__0__anchor__out = cst_27_out1_valid;
	assign cst_27_out1_ready = cst_27__MC_x__ready__0__anchor__in;
	assign cst_27__MC_x__ready__0__anchor__out = MC_x_in2_ready;
	assign MC_w_clk = clk;
	assign MC_w_rst = rst;
	assign w_ce0 = w_we0;
	assign load_80_in1_data = MC_w__load_80__data__0__anchor__in;
	assign MC_w__load_80__data__0__anchor__out = MC_w_out1_data;
	assign load_80_in1_valid = MC_w__load_80__valid__0__anchor__in;
	assign MC_w__load_80__valid__0__anchor__out = MC_w_out1_valid;
	assign MC_w_out1_ready = MC_w__load_80__ready__0__anchor__in;
	assign MC_w__load_80__ready__0__anchor__out = load_80_in1_ready;
	assign end_0_in9_data = MC_w__end_0__data__0__anchor__in;
	assign MC_w__end_0__data__0__anchor__out = MC_w_out2_data;
	assign end_0_in9_valid = MC_w__end_0__valid__0__anchor__in;
	assign MC_w__end_0__valid__0__anchor__out = MC_w_out2_valid;
	assign MC_w_out2_ready = MC_w__end_0__ready__0__anchor__in;
	assign MC_w__end_0__ready__0__anchor__out = end_0_in9_ready;
	assign cst_28_clk = clk;
	assign cst_28_rst = rst;
	assign MC_w_in1_data = cst_28__MC_w__data__0__anchor__in;
	assign cst_28__MC_w__data__0__anchor__out = cst_28_out1_data;
	assign MC_w_in1_valid = cst_28__MC_w__valid__0__anchor__in;
	assign cst_28__MC_w__valid__0__anchor__out = cst_28_out1_valid;
	assign cst_28_out1_ready = cst_28__MC_w__ready__0__anchor__in;
	assign cst_28__MC_w__ready__0__anchor__out = MC_w_in1_ready;
	assign end_0_clk = clk;
	assign end_0_rst = rst;
	assign end_out = end_0_out1_data;
	assign end_0_out1_ready = end_ready;
	assign end_valid = end_0_out1_valid;
	assign start_0_clk = clk;
	assign start_0_rst = rst;
	assign start_0_in1_data = start_in;
	assign start_0_in1_valid = start_valid;
	assign start_ready = start_0_in1_ready;
	assign forkC_44_in1_data = start_0__forkC_44__data__0__anchor__in;
	assign start_0__forkC_44__data__0__anchor__out = start_0_out1_data;
	assign forkC_44_in1_valid = start_0__forkC_44__valid__0__anchor__in;
	assign start_0__forkC_44__valid__0__anchor__out = start_0_out1_valid;
	assign start_0_out1_ready = start_0__forkC_44__ready__0__anchor__in;
	assign start_0__forkC_44__ready__0__anchor__out = forkC_44_in1_ready;
	assign forkC_44_clk = clk;
	assign forkC_44_rst = rst;
	assign cst_0_in1_data = forkC_44__cst_0__data__0__anchor__in;
	assign forkC_44__cst_0__data__0__anchor__out = forkC_44_out1_data;
	assign cst_0_in1_valid = forkC_44__cst_0__valid__0__anchor__in;
	assign forkC_44__cst_0__valid__0__anchor__out = forkC_44_out1_valid;
	assign forkC_44_out1_ready = forkC_44__cst_0__ready__0__anchor__in;
	assign forkC_44__cst_0__ready__0__anchor__out = cst_0_in1_ready;
	assign branchC_46_in1_data = forkC_44__branchC_46__data__0__anchor__in;
	assign forkC_44__branchC_46__data__0__anchor__out = forkC_44_out2_data;
	assign branchC_46_in1_valid = forkC_44__branchC_46__valid__0__anchor__in;
	assign forkC_44__branchC_46__valid__0__anchor__out = forkC_44_out2_valid;
	assign forkC_44_out2_ready = forkC_44__branchC_46__ready__0__anchor__in;
	assign forkC_44__branchC_46__ready__0__anchor__out = branchC_46_in1_ready;
	assign brCst_block1_in1_data = forkC_44__brCst_block1__data__0__anchor__in;
	assign forkC_44__brCst_block1__data__0__anchor__out = forkC_44_out3_data;
	assign brCst_block1_in1_valid = forkC_44__brCst_block1__valid__0__anchor__in;
	assign forkC_44__brCst_block1__valid__0__anchor__out = forkC_44_out3_valid;
	assign forkC_44_out3_ready = forkC_44__brCst_block1__ready__0__anchor__in;
	assign forkC_44__brCst_block1__ready__0__anchor__out = brCst_block1_in1_ready;
	assign branchC_46_clk = clk;
	assign branchC_46_rst = rst;
	assign phiC_28_in1_data = branchC_46__phiC_28__data__0__anchor__in;
	assign branchC_46__phiC_28__data__0__anchor__out = branchC_46_out1_data;
	assign phiC_28_in1_valid = branchC_46__phiC_28__valid__0__anchor__in;
	assign branchC_46__phiC_28__valid__0__anchor__out = branchC_46_out1_valid;
	assign branchC_46_out1_ready = branchC_46__phiC_28__ready__0__anchor__in;
	assign branchC_46__phiC_28__ready__0__anchor__out = phiC_28_in1_ready;
	assign sink_32_in1_data = branchC_46__sink_32__data__0__anchor__in;
	assign branchC_46__sink_32__data__0__anchor__out = branchC_46_out2_data;
	assign sink_32_in1_valid = branchC_46__sink_32__valid__0__anchor__in;
	assign branchC_46__sink_32__valid__0__anchor__out = branchC_46_out2_valid;
	assign branchC_46_out2_ready = branchC_46__sink_32__ready__0__anchor__in;
	assign branchC_46__sink_32__ready__0__anchor__out = sink_32_in1_ready;
	assign phiC_28_clk = clk;
	assign phiC_28_rst = rst;
	assign forkC_45_in1_data = phiC_28__forkC_45__data__0__anchor__in;
	assign phiC_28__forkC_45__data__0__anchor__out = phiC_28_out1_data;
	assign forkC_45_in1_valid = phiC_28__forkC_45__valid__0__anchor__in;
	assign phiC_28__forkC_45__valid__0__anchor__out = phiC_28_out1_valid;
	assign phiC_28_out1_ready = phiC_28__forkC_45__ready__0__anchor__in;
	assign phiC_28__forkC_45__ready__0__anchor__out = forkC_45_in1_ready;
	assign phi_1_in1_data = phiC_28__phi_1__data__0__anchor__in;
	assign phiC_28__phi_1__data__0__anchor__out = phiC_28_out2_data;
	assign phi_1_in1_valid = phiC_28__phi_1__valid__0__anchor__in;
	assign phiC_28__phi_1__valid__0__anchor__out = phiC_28_out2_valid;
	assign phiC_28_out2_ready = phiC_28__phi_1__ready__0__anchor__in;
	assign phiC_28__phi_1__ready__0__anchor__out = phi_1_in1_ready;
	assign forkC_45_clk = clk;
	assign forkC_45_rst = rst;
	assign cst_1_in1_data = forkC_45__cst_1__data__0__anchor__in;
	assign forkC_45__cst_1__data__0__anchor__out = forkC_45_out1_data;
	assign cst_1_in1_valid = forkC_45__cst_1__valid__0__anchor__in;
	assign forkC_45__cst_1__valid__0__anchor__out = forkC_45_out1_valid;
	assign forkC_45_out1_ready = forkC_45__cst_1__ready__0__anchor__in;
	assign forkC_45__cst_1__ready__0__anchor__out = cst_1_in1_ready;
	assign branchC_47_in1_data = forkC_45__branchC_47__data__0__anchor__in;
	assign forkC_45__branchC_47__data__0__anchor__out = forkC_45_out2_data;
	assign branchC_47_in1_valid = forkC_45__branchC_47__valid__0__anchor__in;
	assign forkC_45__branchC_47__valid__0__anchor__out = forkC_45_out2_valid;
	assign forkC_45_out2_ready = forkC_45__branchC_47__ready__0__anchor__in;
	assign forkC_45__branchC_47__ready__0__anchor__out = branchC_47_in1_ready;
	assign brCst_block2_in1_data = forkC_45__brCst_block2__data__0__anchor__in;
	assign forkC_45__brCst_block2__data__0__anchor__out = forkC_45_out3_data;
	assign brCst_block2_in1_valid = forkC_45__brCst_block2__valid__0__anchor__in;
	assign forkC_45__brCst_block2__valid__0__anchor__out = forkC_45_out3_valid;
	assign forkC_45_out3_ready = forkC_45__brCst_block2__ready__0__anchor__in;
	assign forkC_45__brCst_block2__ready__0__anchor__out = brCst_block2_in1_ready;
	assign branchC_47_clk = clk;
	assign branchC_47_rst = rst;
	assign phiC_29_in1_data = branchC_47__phiC_29__data__0__anchor__in;
	assign branchC_47__phiC_29__data__0__anchor__out = branchC_47_out1_data;
	assign phiC_29_in1_valid = branchC_47__phiC_29__valid__0__anchor__in;
	assign branchC_47__phiC_29__valid__0__anchor__out = branchC_47_out1_valid;
	assign branchC_47_out1_ready = branchC_47__phiC_29__ready__0__anchor__in;
	assign branchC_47__phiC_29__ready__0__anchor__out = phiC_29_in1_ready;
	assign sink_33_in1_data = branchC_47__sink_33__data__0__anchor__in;
	assign branchC_47__sink_33__data__0__anchor__out = branchC_47_out2_data;
	assign sink_33_in1_valid = branchC_47__sink_33__valid__0__anchor__in;
	assign branchC_47__sink_33__valid__0__anchor__out = branchC_47_out2_valid;
	assign branchC_47_out2_ready = branchC_47__sink_33__ready__0__anchor__in;
	assign branchC_47__sink_33__ready__0__anchor__out = sink_33_in1_ready;
	assign phiC_29_clk = clk;
	assign phiC_29_rst = rst;
	assign forkC_46_in1_data = phiC_29__forkC_46__data__0__anchor__in;
	assign phiC_29__forkC_46__data__0__anchor__out = phiC_29_out1_data;
	assign forkC_46_in1_valid = phiC_29__forkC_46__valid__0__anchor__in;
	assign phiC_29__forkC_46__valid__0__anchor__out = phiC_29_out1_valid;
	assign phiC_29_out1_ready = phiC_29__forkC_46__ready__0__anchor__in;
	assign phiC_29__forkC_46__ready__0__anchor__out = forkC_46_in1_ready;
	assign phi_3_in1_data = phiC_29__phi_3__data__0__anchor__in;
	assign phiC_29__phi_3__data__0__anchor__out = phiC_29_out2_data;
	assign phi_3_in1_valid = phiC_29__phi_3__valid__0__anchor__in;
	assign phiC_29__phi_3__valid__0__anchor__out = phiC_29_out2_valid;
	assign phiC_29_out2_ready = phiC_29__phi_3__ready__0__anchor__in;
	assign phiC_29__phi_3__ready__0__anchor__out = phi_3_in1_ready;
	assign forkC_46_clk = clk;
	assign forkC_46_rst = rst;
	assign cst_25_in1_data = forkC_46__cst_25__data__0__anchor__in;
	assign forkC_46__cst_25__data__0__anchor__out = forkC_46_out1_data;
	assign cst_25_in1_valid = forkC_46__cst_25__valid__0__anchor__in;
	assign forkC_46__cst_25__valid__0__anchor__out = forkC_46_out1_valid;
	assign forkC_46_out1_ready = forkC_46__cst_25__ready__0__anchor__in;
	assign forkC_46__cst_25__ready__0__anchor__out = cst_25_in1_ready;
	assign branchC_48_in1_data = forkC_46__branchC_48__data__0__anchor__in;
	assign forkC_46__branchC_48__data__0__anchor__out = forkC_46_out2_data;
	assign branchC_48_in1_valid = forkC_46__branchC_48__valid__0__anchor__in;
	assign forkC_46__branchC_48__valid__0__anchor__out = forkC_46_out2_valid;
	assign forkC_46_out2_ready = forkC_46__branchC_48__ready__0__anchor__in;
	assign forkC_46__branchC_48__ready__0__anchor__out = branchC_48_in1_ready;
	assign branchC_48_clk = clk;
	assign branchC_48_rst = rst;
	assign Buffer_20_in1_data = branchC_48__Buffer_20__data__0__anchor__in;
	assign branchC_48__Buffer_20__data__0__anchor__out = branchC_48_out1_data;
	assign Buffer_20_in1_valid = branchC_48__Buffer_20__valid__0__anchor__in;
	assign branchC_48__Buffer_20__valid__0__anchor__out = branchC_48_out1_valid;
	assign branchC_48_out1_ready = branchC_48__Buffer_20__ready__0__anchor__in;
	assign branchC_48__Buffer_20__ready__0__anchor__out = Buffer_20_in1_ready;
	assign phiC_30_in1_data = branchC_48__phiC_30__data__0__anchor__in;
	assign branchC_48__phiC_30__data__0__anchor__out = branchC_48_out2_data;
	assign phiC_30_in1_valid = branchC_48__phiC_30__valid__0__anchor__in;
	assign branchC_48__phiC_30__valid__0__anchor__out = branchC_48_out2_valid;
	assign branchC_48_out2_ready = branchC_48__phiC_30__ready__0__anchor__in;
	assign branchC_48__phiC_30__ready__0__anchor__out = phiC_30_in1_ready;
	assign phiC_30_clk = clk;
	assign phiC_30_rst = rst;
	assign branchC_49_in1_data = phiC_30__branchC_49__data__0__anchor__in;
	assign phiC_30__branchC_49__data__0__anchor__out = phiC_30_out1_data;
	assign branchC_49_in1_valid = phiC_30__branchC_49__valid__0__anchor__in;
	assign phiC_30__branchC_49__valid__0__anchor__out = phiC_30_out1_valid;
	assign phiC_30_out1_ready = phiC_30__branchC_49__ready__0__anchor__in;
	assign phiC_30__branchC_49__ready__0__anchor__out = branchC_49_in1_ready;
	assign branchC_49_clk = clk;
	assign branchC_49_rst = rst;
	assign Buffer_16_in1_data = branchC_49__Buffer_16__data__0__anchor__in;
	assign branchC_49__Buffer_16__data__0__anchor__out = branchC_49_out1_data;
	assign Buffer_16_in1_valid = branchC_49__Buffer_16__valid__0__anchor__in;
	assign branchC_49__Buffer_16__valid__0__anchor__out = branchC_49_out1_valid;
	assign branchC_49_out1_ready = branchC_49__Buffer_16__ready__0__anchor__in;
	assign branchC_49__Buffer_16__ready__0__anchor__out = Buffer_16_in1_ready;
	assign phiC_31_in1_data = branchC_49__phiC_31__data__0__anchor__in;
	assign branchC_49__phiC_31__data__0__anchor__out = branchC_49_out2_data;
	assign phiC_31_in1_valid = branchC_49__phiC_31__valid__0__anchor__in;
	assign branchC_49__phiC_31__valid__0__anchor__out = branchC_49_out2_valid;
	assign branchC_49_out2_ready = branchC_49__phiC_31__ready__0__anchor__in;
	assign branchC_49__phiC_31__ready__0__anchor__out = phiC_31_in1_ready;
	assign phiC_31_clk = clk;
	assign phiC_31_rst = rst;
	assign forkC_48_in1_data = phiC_31__forkC_48__data__0__anchor__in;
	assign phiC_31__forkC_48__data__0__anchor__out = phiC_31_out1_data;
	assign forkC_48_in1_valid = phiC_31__forkC_48__valid__0__anchor__in;
	assign phiC_31__forkC_48__valid__0__anchor__out = phiC_31_out1_valid;
	assign phiC_31_out1_ready = phiC_31__forkC_48__ready__0__anchor__in;
	assign phiC_31__forkC_48__ready__0__anchor__out = forkC_48_in1_ready;
	assign forkC_48_clk = clk;
	assign forkC_48_rst = rst;
	assign cst_8_in1_data = forkC_48__cst_8__data__0__anchor__in;
	assign forkC_48__cst_8__data__0__anchor__out = forkC_48_out1_data;
	assign cst_8_in1_valid = forkC_48__cst_8__valid__0__anchor__in;
	assign forkC_48__cst_8__valid__0__anchor__out = forkC_48_out1_valid;
	assign forkC_48_out1_ready = forkC_48__cst_8__ready__0__anchor__in;
	assign forkC_48__cst_8__ready__0__anchor__out = cst_8_in1_ready;
	assign branchC_50_in1_data = forkC_48__branchC_50__data__0__anchor__in;
	assign forkC_48__branchC_50__data__0__anchor__out = forkC_48_out2_data;
	assign branchC_50_in1_valid = forkC_48__branchC_50__valid__0__anchor__in;
	assign forkC_48__branchC_50__valid__0__anchor__out = forkC_48_out2_valid;
	assign forkC_48_out2_ready = forkC_48__branchC_50__ready__0__anchor__in;
	assign forkC_48__branchC_50__ready__0__anchor__out = branchC_50_in1_ready;
	assign brCst_block5_in1_data = forkC_48__brCst_block5__data__0__anchor__in;
	assign forkC_48__brCst_block5__data__0__anchor__out = forkC_48_out3_data;
	assign brCst_block5_in1_valid = forkC_48__brCst_block5__valid__0__anchor__in;
	assign forkC_48__brCst_block5__valid__0__anchor__out = forkC_48_out3_valid;
	assign forkC_48_out3_ready = forkC_48__brCst_block5__ready__0__anchor__in;
	assign forkC_48__brCst_block5__ready__0__anchor__out = brCst_block5_in1_ready;
	assign branchC_50_clk = clk;
	assign branchC_50_rst = rst;
	assign phiC_32_in1_data = branchC_50__phiC_32__data__0__anchor__in;
	assign branchC_50__phiC_32__data__0__anchor__out = branchC_50_out1_data;
	assign phiC_32_in1_valid = branchC_50__phiC_32__valid__0__anchor__in;
	assign branchC_50__phiC_32__valid__0__anchor__out = branchC_50_out1_valid;
	assign branchC_50_out1_ready = branchC_50__phiC_32__ready__0__anchor__in;
	assign branchC_50__phiC_32__ready__0__anchor__out = phiC_32_in1_ready;
	assign sink_34_in1_data = branchC_50__sink_34__data__0__anchor__in;
	assign branchC_50__sink_34__data__0__anchor__out = branchC_50_out2_data;
	assign sink_34_in1_valid = branchC_50__sink_34__valid__0__anchor__in;
	assign branchC_50__sink_34__valid__0__anchor__out = branchC_50_out2_valid;
	assign branchC_50_out2_ready = branchC_50__sink_34__ready__0__anchor__in;
	assign branchC_50__sink_34__ready__0__anchor__out = sink_34_in1_ready;
	assign phiC_32_clk = clk;
	assign phiC_32_rst = rst;
	assign forkC_49_in1_data = phiC_32__forkC_49__data__0__anchor__in;
	assign phiC_32__forkC_49__data__0__anchor__out = phiC_32_out1_data;
	assign forkC_49_in1_valid = phiC_32__forkC_49__valid__0__anchor__in;
	assign phiC_32__forkC_49__valid__0__anchor__out = phiC_32_out1_valid;
	assign phiC_32_out1_ready = phiC_32__forkC_49__ready__0__anchor__in;
	assign phiC_32__forkC_49__ready__0__anchor__out = forkC_49_in1_ready;
	assign phi_36_in1_data = phiC_32__phi_36__data__0__anchor__in;
	assign phiC_32__phi_36__data__0__anchor__out = phiC_32_out2_data;
	assign phi_36_in1_valid = phiC_32__phi_36__valid__0__anchor__in;
	assign phiC_32__phi_36__valid__0__anchor__out = phiC_32_out2_valid;
	assign phiC_32_out2_ready = phiC_32__phi_36__ready__0__anchor__in;
	assign phiC_32__phi_36__ready__0__anchor__out = phi_36_in1_ready;
	assign forkC_49_clk = clk;
	assign forkC_49_rst = rst;
	assign cst_9_in1_data = forkC_49__cst_9__data__0__anchor__in;
	assign forkC_49__cst_9__data__0__anchor__out = forkC_49_out1_data;
	assign cst_9_in1_valid = forkC_49__cst_9__valid__0__anchor__in;
	assign forkC_49__cst_9__valid__0__anchor__out = forkC_49_out1_valid;
	assign forkC_49_out1_ready = forkC_49__cst_9__ready__0__anchor__in;
	assign forkC_49__cst_9__ready__0__anchor__out = cst_9_in1_ready;
	assign branchC_51_in1_data = forkC_49__branchC_51__data__0__anchor__in;
	assign forkC_49__branchC_51__data__0__anchor__out = forkC_49_out2_data;
	assign branchC_51_in1_valid = forkC_49__branchC_51__valid__0__anchor__in;
	assign forkC_49__branchC_51__valid__0__anchor__out = forkC_49_out2_valid;
	assign forkC_49_out2_ready = forkC_49__branchC_51__ready__0__anchor__in;
	assign forkC_49__branchC_51__ready__0__anchor__out = branchC_51_in1_ready;
	assign brCst_block6_in1_data = forkC_49__brCst_block6__data__0__anchor__in;
	assign forkC_49__brCst_block6__data__0__anchor__out = forkC_49_out3_data;
	assign brCst_block6_in1_valid = forkC_49__brCst_block6__valid__0__anchor__in;
	assign forkC_49__brCst_block6__valid__0__anchor__out = forkC_49_out3_valid;
	assign forkC_49_out3_ready = forkC_49__brCst_block6__ready__0__anchor__in;
	assign forkC_49__brCst_block6__ready__0__anchor__out = brCst_block6_in1_ready;
	assign branchC_51_clk = clk;
	assign branchC_51_rst = rst;
	assign phiC_33_in1_data = branchC_51__phiC_33__data__0__anchor__in;
	assign branchC_51__phiC_33__data__0__anchor__out = branchC_51_out1_data;
	assign phiC_33_in1_valid = branchC_51__phiC_33__valid__0__anchor__in;
	assign branchC_51__phiC_33__valid__0__anchor__out = branchC_51_out1_valid;
	assign branchC_51_out1_ready = branchC_51__phiC_33__ready__0__anchor__in;
	assign branchC_51__phiC_33__ready__0__anchor__out = phiC_33_in1_ready;
	assign sink_35_in1_data = branchC_51__sink_35__data__0__anchor__in;
	assign branchC_51__sink_35__data__0__anchor__out = branchC_51_out2_data;
	assign sink_35_in1_valid = branchC_51__sink_35__valid__0__anchor__in;
	assign branchC_51__sink_35__valid__0__anchor__out = branchC_51_out2_valid;
	assign branchC_51_out2_ready = branchC_51__sink_35__ready__0__anchor__in;
	assign branchC_51__sink_35__ready__0__anchor__out = sink_35_in1_ready;
	assign phiC_33_clk = clk;
	assign phiC_33_rst = rst;
	assign branchC_52_in1_data = phiC_33__branchC_52__data__0__anchor__in;
	assign phiC_33__branchC_52__data__0__anchor__out = phiC_33_out1_data;
	assign branchC_52_in1_valid = phiC_33__branchC_52__valid__0__anchor__in;
	assign phiC_33__branchC_52__valid__0__anchor__out = phiC_33_out1_valid;
	assign phiC_33_out1_ready = phiC_33__branchC_52__ready__0__anchor__in;
	assign phiC_33__branchC_52__ready__0__anchor__out = branchC_52_in1_ready;
	assign fork_62_in1_data = phiC_33__fork_62__data__0__anchor__in;
	assign phiC_33__fork_62__data__0__anchor__out = phiC_33_out2_data;
	assign fork_62_in1_valid = phiC_33__fork_62__valid__0__anchor__in;
	assign phiC_33__fork_62__valid__0__anchor__out = phiC_33_out2_valid;
	assign phiC_33_out2_ready = phiC_33__fork_62__ready__0__anchor__in;
	assign phiC_33__fork_62__ready__0__anchor__out = fork_62_in1_ready;
	assign branchC_52_clk = clk;
	assign branchC_52_rst = rst;
	assign Buffer_21_in1_data = branchC_52__Buffer_21__data__0__anchor__in;
	assign branchC_52__Buffer_21__data__0__anchor__out = branchC_52_out1_data;
	assign Buffer_21_in1_valid = branchC_52__Buffer_21__valid__0__anchor__in;
	assign branchC_52__Buffer_21__valid__0__anchor__out = branchC_52_out1_valid;
	assign branchC_52_out1_ready = branchC_52__Buffer_21__ready__0__anchor__in;
	assign branchC_52__Buffer_21__ready__0__anchor__out = Buffer_21_in1_ready;
	assign phiC_34_in1_data = branchC_52__phiC_34__data__0__anchor__in;
	assign branchC_52__phiC_34__data__0__anchor__out = branchC_52_out2_data;
	assign phiC_34_in1_valid = branchC_52__phiC_34__valid__0__anchor__in;
	assign branchC_52__phiC_34__valid__0__anchor__out = branchC_52_out2_valid;
	assign branchC_52_out2_ready = branchC_52__phiC_34__ready__0__anchor__in;
	assign branchC_52__phiC_34__ready__0__anchor__out = phiC_34_in1_ready;
	assign phiC_34_clk = clk;
	assign phiC_34_rst = rst;
	assign forkC_51_in1_data = phiC_34__forkC_51__data__0__anchor__in;
	assign phiC_34__forkC_51__data__0__anchor__out = phiC_34_out1_data;
	assign forkC_51_in1_valid = phiC_34__forkC_51__valid__0__anchor__in;
	assign phiC_34__forkC_51__valid__0__anchor__out = phiC_34_out1_valid;
	assign phiC_34_out1_ready = phiC_34__forkC_51__ready__0__anchor__in;
	assign phiC_34__forkC_51__ready__0__anchor__out = forkC_51_in1_ready;
	assign forkC_51_clk = clk;
	assign forkC_51_rst = rst;
	assign cst_26_in1_data = forkC_51__cst_26__data__0__anchor__in;
	assign forkC_51__cst_26__data__0__anchor__out = forkC_51_out1_data;
	assign cst_26_in1_valid = forkC_51__cst_26__valid__0__anchor__in;
	assign forkC_51__cst_26__valid__0__anchor__out = forkC_51_out1_valid;
	assign forkC_51_out1_ready = forkC_51__cst_26__ready__0__anchor__in;
	assign forkC_51__cst_26__ready__0__anchor__out = cst_26_in1_ready;
	assign branchC_53_in1_data = forkC_51__branchC_53__data__0__anchor__in;
	assign forkC_51__branchC_53__data__0__anchor__out = forkC_51_out2_data;
	assign branchC_53_in1_valid = forkC_51__branchC_53__valid__0__anchor__in;
	assign forkC_51__branchC_53__valid__0__anchor__out = forkC_51_out2_valid;
	assign forkC_51_out2_ready = forkC_51__branchC_53__ready__0__anchor__in;
	assign forkC_51__branchC_53__ready__0__anchor__out = branchC_53_in1_ready;
	assign branchC_53_clk = clk;
	assign branchC_53_rst = rst;
	assign Buffer_27_in1_data = branchC_53__Buffer_27__data__0__anchor__in;
	assign branchC_53__Buffer_27__data__0__anchor__out = branchC_53_out1_data;
	assign Buffer_27_in1_valid = branchC_53__Buffer_27__valid__0__anchor__in;
	assign branchC_53__Buffer_27__valid__0__anchor__out = branchC_53_out1_valid;
	assign branchC_53_out1_ready = branchC_53__Buffer_27__ready__0__anchor__in;
	assign branchC_53__Buffer_27__ready__0__anchor__out = Buffer_27_in1_ready;
	assign phiC_35_in1_data = branchC_53__phiC_35__data__0__anchor__in;
	assign branchC_53__phiC_35__data__0__anchor__out = branchC_53_out2_data;
	assign phiC_35_in1_valid = branchC_53__phiC_35__valid__0__anchor__in;
	assign branchC_53__phiC_35__valid__0__anchor__out = branchC_53_out2_valid;
	assign branchC_53_out2_ready = branchC_53__phiC_35__ready__0__anchor__in;
	assign branchC_53__phiC_35__ready__0__anchor__out = phiC_35_in1_ready;
	assign phiC_35_clk = clk;
	assign phiC_35_rst = rst;
	assign forkC_52_in1_data = phiC_35__forkC_52__data__0__anchor__in;
	assign phiC_35__forkC_52__data__0__anchor__out = phiC_35_out1_data;
	assign forkC_52_in1_valid = phiC_35__forkC_52__valid__0__anchor__in;
	assign phiC_35__forkC_52__valid__0__anchor__out = phiC_35_out1_valid;
	assign phiC_35_out1_ready = phiC_35__forkC_52__ready__0__anchor__in;
	assign phiC_35__forkC_52__ready__0__anchor__out = forkC_52_in1_ready;
	assign forkC_52_clk = clk;
	assign forkC_52_rst = rst;
	assign cst_15_in1_data = forkC_52__cst_15__data__0__anchor__in;
	assign forkC_52__cst_15__data__0__anchor__out = forkC_52_out1_data;
	assign cst_15_in1_valid = forkC_52__cst_15__valid__0__anchor__in;
	assign forkC_52__cst_15__valid__0__anchor__out = forkC_52_out1_valid;
	assign forkC_52_out1_ready = forkC_52__cst_15__ready__0__anchor__in;
	assign forkC_52__cst_15__ready__0__anchor__out = cst_15_in1_ready;
	assign branchC_54_in1_data = forkC_52__branchC_54__data__0__anchor__in;
	assign forkC_52__branchC_54__data__0__anchor__out = forkC_52_out2_data;
	assign branchC_54_in1_valid = forkC_52__branchC_54__valid__0__anchor__in;
	assign forkC_52__branchC_54__valid__0__anchor__out = forkC_52_out2_valid;
	assign forkC_52_out2_ready = forkC_52__branchC_54__ready__0__anchor__in;
	assign forkC_52__branchC_54__ready__0__anchor__out = branchC_54_in1_ready;
	assign brCst_block9_in1_data = forkC_52__brCst_block9__data__0__anchor__in;
	assign forkC_52__brCst_block9__data__0__anchor__out = forkC_52_out3_data;
	assign brCst_block9_in1_valid = forkC_52__brCst_block9__valid__0__anchor__in;
	assign forkC_52__brCst_block9__valid__0__anchor__out = forkC_52_out3_valid;
	assign forkC_52_out3_ready = forkC_52__brCst_block9__ready__0__anchor__in;
	assign forkC_52__brCst_block9__ready__0__anchor__out = brCst_block9_in1_ready;
	assign branchC_54_clk = clk;
	assign branchC_54_rst = rst;
	assign phiC_36_in1_data = branchC_54__phiC_36__data__0__anchor__in;
	assign branchC_54__phiC_36__data__0__anchor__out = branchC_54_out1_data;
	assign phiC_36_in1_valid = branchC_54__phiC_36__valid__0__anchor__in;
	assign branchC_54__phiC_36__valid__0__anchor__out = branchC_54_out1_valid;
	assign branchC_54_out1_ready = branchC_54__phiC_36__ready__0__anchor__in;
	assign branchC_54__phiC_36__ready__0__anchor__out = phiC_36_in1_ready;
	assign sink_36_in1_data = branchC_54__sink_36__data__0__anchor__in;
	assign branchC_54__sink_36__data__0__anchor__out = branchC_54_out2_data;
	assign sink_36_in1_valid = branchC_54__sink_36__valid__0__anchor__in;
	assign branchC_54__sink_36__valid__0__anchor__out = branchC_54_out2_valid;
	assign branchC_54_out2_ready = branchC_54__sink_36__ready__0__anchor__in;
	assign branchC_54__sink_36__ready__0__anchor__out = sink_36_in1_ready;
	assign phiC_36_clk = clk;
	assign phiC_36_rst = rst;
	assign forkC_53_in1_data = phiC_36__forkC_53__data__0__anchor__in;
	assign phiC_36__forkC_53__data__0__anchor__out = phiC_36_out1_data;
	assign forkC_53_in1_valid = phiC_36__forkC_53__valid__0__anchor__in;
	assign phiC_36__forkC_53__valid__0__anchor__out = phiC_36_out1_valid;
	assign phiC_36_out1_ready = phiC_36__forkC_53__ready__0__anchor__in;
	assign phiC_36__forkC_53__ready__0__anchor__out = forkC_53_in1_ready;
	assign phi_63_in1_data = phiC_36__phi_63__data__0__anchor__in;
	assign phiC_36__phi_63__data__0__anchor__out = phiC_36_out2_data;
	assign phi_63_in1_valid = phiC_36__phi_63__valid__0__anchor__in;
	assign phiC_36__phi_63__valid__0__anchor__out = phiC_36_out2_valid;
	assign phiC_36_out2_ready = phiC_36__phi_63__ready__0__anchor__in;
	assign phiC_36__phi_63__ready__0__anchor__out = phi_63_in1_ready;
	assign forkC_53_clk = clk;
	assign forkC_53_rst = rst;
	assign cst_27_in1_data = forkC_53__cst_27__data__0__anchor__in;
	assign forkC_53__cst_27__data__0__anchor__out = forkC_53_out1_data;
	assign cst_27_in1_valid = forkC_53__cst_27__valid__0__anchor__in;
	assign forkC_53__cst_27__valid__0__anchor__out = forkC_53_out1_valid;
	assign forkC_53_out1_ready = forkC_53__cst_27__ready__0__anchor__in;
	assign forkC_53__cst_27__ready__0__anchor__out = cst_27_in1_ready;
	assign branchC_55_in1_data = forkC_53__branchC_55__data__0__anchor__in;
	assign forkC_53__branchC_55__data__0__anchor__out = forkC_53_out2_data;
	assign branchC_55_in1_valid = forkC_53__branchC_55__valid__0__anchor__in;
	assign forkC_53__branchC_55__valid__0__anchor__out = forkC_53_out2_valid;
	assign forkC_53_out2_ready = forkC_53__branchC_55__ready__0__anchor__in;
	assign forkC_53__branchC_55__ready__0__anchor__out = branchC_55_in1_ready;
	assign branchC_55_clk = clk;
	assign branchC_55_rst = rst;
	assign Buffer_7_in1_data = branchC_55__Buffer_7__data__0__anchor__in;
	assign branchC_55__Buffer_7__data__0__anchor__out = branchC_55_out1_data;
	assign Buffer_7_in1_valid = branchC_55__Buffer_7__valid__0__anchor__in;
	assign branchC_55__Buffer_7__valid__0__anchor__out = branchC_55_out1_valid;
	assign branchC_55_out1_ready = branchC_55__Buffer_7__ready__0__anchor__in;
	assign branchC_55__Buffer_7__ready__0__anchor__out = Buffer_7_in1_ready;
	assign phiC_37_in1_data = branchC_55__phiC_37__data__0__anchor__in;
	assign branchC_55__phiC_37__data__0__anchor__out = branchC_55_out2_data;
	assign phiC_37_in1_valid = branchC_55__phiC_37__valid__0__anchor__in;
	assign branchC_55__phiC_37__valid__0__anchor__out = branchC_55_out2_valid;
	assign branchC_55_out2_ready = branchC_55__phiC_37__ready__0__anchor__in;
	assign branchC_55__phiC_37__ready__0__anchor__out = phiC_37_in1_ready;
	assign phiC_37_clk = clk;
	assign phiC_37_rst = rst;
	assign forkC_54_in1_data = phiC_37__forkC_54__data__0__anchor__in;
	assign phiC_37__forkC_54__data__0__anchor__out = phiC_37_out1_data;
	assign forkC_54_in1_valid = phiC_37__forkC_54__valid__0__anchor__in;
	assign phiC_37__forkC_54__valid__0__anchor__out = phiC_37_out1_valid;
	assign phiC_37_out1_ready = phiC_37__forkC_54__ready__0__anchor__in;
	assign phiC_37__forkC_54__ready__0__anchor__out = forkC_54_in1_ready;
	assign forkC_54_clk = clk;
	assign forkC_54_rst = rst;
	assign cst_18_in1_data = forkC_54__cst_18__data__0__anchor__in;
	assign forkC_54__cst_18__data__0__anchor__out = forkC_54_out1_data;
	assign cst_18_in1_valid = forkC_54__cst_18__valid__0__anchor__in;
	assign forkC_54__cst_18__valid__0__anchor__out = forkC_54_out1_valid;
	assign forkC_54_out1_ready = forkC_54__cst_18__ready__0__anchor__in;
	assign forkC_54__cst_18__ready__0__anchor__out = cst_18_in1_ready;
	assign branchC_56_in1_data = forkC_54__branchC_56__data__0__anchor__in;
	assign forkC_54__branchC_56__data__0__anchor__out = forkC_54_out2_data;
	assign branchC_56_in1_valid = forkC_54__branchC_56__valid__0__anchor__in;
	assign forkC_54__branchC_56__valid__0__anchor__out = forkC_54_out2_valid;
	assign forkC_54_out2_ready = forkC_54__branchC_56__ready__0__anchor__in;
	assign forkC_54__branchC_56__ready__0__anchor__out = branchC_56_in1_ready;
	assign brCst_block11_in1_data = forkC_54__brCst_block11__data__0__anchor__in;
	assign forkC_54__brCst_block11__data__0__anchor__out = forkC_54_out3_data;
	assign brCst_block11_in1_valid = forkC_54__brCst_block11__valid__0__anchor__in;
	assign forkC_54__brCst_block11__valid__0__anchor__out = forkC_54_out3_valid;
	assign forkC_54_out3_ready = forkC_54__brCst_block11__ready__0__anchor__in;
	assign forkC_54__brCst_block11__ready__0__anchor__out = brCst_block11_in1_ready;
	assign branchC_56_clk = clk;
	assign branchC_56_rst = rst;
	assign phiC_38_in1_data = branchC_56__phiC_38__data__0__anchor__in;
	assign branchC_56__phiC_38__data__0__anchor__out = branchC_56_out1_data;
	assign phiC_38_in1_valid = branchC_56__phiC_38__valid__0__anchor__in;
	assign branchC_56__phiC_38__valid__0__anchor__out = branchC_56_out1_valid;
	assign branchC_56_out1_ready = branchC_56__phiC_38__ready__0__anchor__in;
	assign branchC_56__phiC_38__ready__0__anchor__out = phiC_38_in1_ready;
	assign sink_37_in1_data = branchC_56__sink_37__data__0__anchor__in;
	assign branchC_56__sink_37__data__0__anchor__out = branchC_56_out2_data;
	assign sink_37_in1_valid = branchC_56__sink_37__valid__0__anchor__in;
	assign branchC_56__sink_37__valid__0__anchor__out = branchC_56_out2_valid;
	assign branchC_56_out2_ready = branchC_56__sink_37__ready__0__anchor__in;
	assign branchC_56__sink_37__ready__0__anchor__out = sink_37_in1_ready;
	assign phiC_38_clk = clk;
	assign phiC_38_rst = rst;
	assign Buffer_30_in1_data = phiC_38__Buffer_30__data__0__anchor__in;
	assign phiC_38__Buffer_30__data__0__anchor__out = phiC_38_out1_data;
	assign Buffer_30_in1_valid = phiC_38__Buffer_30__valid__0__anchor__in;
	assign phiC_38__Buffer_30__valid__0__anchor__out = phiC_38_out1_valid;
	assign phiC_38_out1_ready = phiC_38__Buffer_30__ready__0__anchor__in;
	assign phiC_38__Buffer_30__ready__0__anchor__out = Buffer_30_in1_ready;
	assign phi_77_in1_data = phiC_38__phi_77__data__0__anchor__in;
	assign phiC_38__phi_77__data__0__anchor__out = phiC_38_out2_data;
	assign phi_77_in1_valid = phiC_38__phi_77__valid__0__anchor__in;
	assign phiC_38__phi_77__valid__0__anchor__out = phiC_38_out2_valid;
	assign phiC_38_out2_ready = phiC_38__phi_77__ready__0__anchor__in;
	assign phiC_38__phi_77__ready__0__anchor__out = phi_77_in1_ready;
	assign forkC_55_clk = clk;
	assign forkC_55_rst = rst;
	assign cst_19_in1_data = forkC_55__cst_19__data__0__anchor__in;
	assign forkC_55__cst_19__data__0__anchor__out = forkC_55_out1_data;
	assign cst_19_in1_valid = forkC_55__cst_19__valid__0__anchor__in;
	assign forkC_55__cst_19__valid__0__anchor__out = forkC_55_out1_valid;
	assign forkC_55_out1_ready = forkC_55__cst_19__ready__0__anchor__in;
	assign forkC_55__cst_19__ready__0__anchor__out = cst_19_in1_ready;
	assign branchC_57_in1_data = forkC_55__branchC_57__data__0__anchor__in;
	assign forkC_55__branchC_57__data__0__anchor__out = forkC_55_out2_data;
	assign branchC_57_in1_valid = forkC_55__branchC_57__valid__0__anchor__in;
	assign forkC_55__branchC_57__valid__0__anchor__out = forkC_55_out2_valid;
	assign forkC_55_out2_ready = forkC_55__branchC_57__ready__0__anchor__in;
	assign forkC_55__branchC_57__ready__0__anchor__out = branchC_57_in1_ready;
	assign brCst_block12_in1_data = forkC_55__brCst_block12__data__0__anchor__in;
	assign forkC_55__brCst_block12__data__0__anchor__out = forkC_55_out3_data;
	assign brCst_block12_in1_valid = forkC_55__brCst_block12__valid__0__anchor__in;
	assign forkC_55__brCst_block12__valid__0__anchor__out = forkC_55_out3_valid;
	assign forkC_55_out3_ready = forkC_55__brCst_block12__ready__0__anchor__in;
	assign forkC_55__brCst_block12__ready__0__anchor__out = brCst_block12_in1_ready;
	assign branchC_57_clk = clk;
	assign branchC_57_rst = rst;
	assign phiC_39_in1_data = branchC_57__phiC_39__data__0__anchor__in;
	assign branchC_57__phiC_39__data__0__anchor__out = branchC_57_out1_data;
	assign phiC_39_in1_valid = branchC_57__phiC_39__valid__0__anchor__in;
	assign branchC_57__phiC_39__valid__0__anchor__out = branchC_57_out1_valid;
	assign branchC_57_out1_ready = branchC_57__phiC_39__ready__0__anchor__in;
	assign branchC_57__phiC_39__ready__0__anchor__out = phiC_39_in1_ready;
	assign sink_38_in1_data = branchC_57__sink_38__data__0__anchor__in;
	assign branchC_57__sink_38__data__0__anchor__out = branchC_57_out2_data;
	assign sink_38_in1_valid = branchC_57__sink_38__valid__0__anchor__in;
	assign branchC_57__sink_38__valid__0__anchor__out = branchC_57_out2_valid;
	assign branchC_57_out2_ready = branchC_57__sink_38__ready__0__anchor__in;
	assign branchC_57__sink_38__ready__0__anchor__out = sink_38_in1_ready;
	assign phiC_39_clk = clk;
	assign phiC_39_rst = rst;
	assign branchC_58_in1_data = phiC_39__branchC_58__data__0__anchor__in;
	assign phiC_39__branchC_58__data__0__anchor__out = phiC_39_out1_data;
	assign branchC_58_in1_valid = phiC_39__branchC_58__valid__0__anchor__in;
	assign phiC_39__branchC_58__valid__0__anchor__out = phiC_39_out1_valid;
	assign phiC_39_out1_ready = phiC_39__branchC_58__ready__0__anchor__in;
	assign phiC_39__branchC_58__ready__0__anchor__out = branchC_58_in1_ready;
	assign fork_65_in1_data = phiC_39__fork_65__data__0__anchor__in;
	assign phiC_39__fork_65__data__0__anchor__out = phiC_39_out2_data;
	assign fork_65_in1_valid = phiC_39__fork_65__valid__0__anchor__in;
	assign phiC_39__fork_65__valid__0__anchor__out = phiC_39_out2_valid;
	assign phiC_39_out2_ready = phiC_39__fork_65__ready__0__anchor__in;
	assign phiC_39__fork_65__ready__0__anchor__out = fork_65_in1_ready;
	assign branchC_58_clk = clk;
	assign branchC_58_rst = rst;
	assign Buffer_2_in1_data = branchC_58__Buffer_2__data__0__anchor__in;
	assign branchC_58__Buffer_2__data__0__anchor__out = branchC_58_out1_data;
	assign Buffer_2_in1_valid = branchC_58__Buffer_2__valid__0__anchor__in;
	assign branchC_58__Buffer_2__valid__0__anchor__out = branchC_58_out1_valid;
	assign branchC_58_out1_ready = branchC_58__Buffer_2__ready__0__anchor__in;
	assign branchC_58__Buffer_2__ready__0__anchor__out = Buffer_2_in1_ready;
	assign phiC_40_in1_data = branchC_58__phiC_40__data__0__anchor__in;
	assign branchC_58__phiC_40__data__0__anchor__out = branchC_58_out2_data;
	assign phiC_40_in1_valid = branchC_58__phiC_40__valid__0__anchor__in;
	assign branchC_58__phiC_40__valid__0__anchor__out = branchC_58_out2_valid;
	assign branchC_58_out2_ready = branchC_58__phiC_40__ready__0__anchor__in;
	assign branchC_58__phiC_40__ready__0__anchor__out = phiC_40_in1_ready;
	assign phiC_40_clk = clk;
	assign phiC_40_rst = rst;
	assign forkC_57_in1_data = phiC_40__forkC_57__data__0__anchor__in;
	assign phiC_40__forkC_57__data__0__anchor__out = phiC_40_out1_data;
	assign forkC_57_in1_valid = phiC_40__forkC_57__valid__0__anchor__in;
	assign phiC_40__forkC_57__valid__0__anchor__out = phiC_40_out1_valid;
	assign phiC_40_out1_ready = phiC_40__forkC_57__ready__0__anchor__in;
	assign phiC_40__forkC_57__ready__0__anchor__out = forkC_57_in1_ready;
	assign forkC_57_clk = clk;
	assign forkC_57_rst = rst;
	assign cst_28_in1_data = forkC_57__cst_28__data__0__anchor__in;
	assign forkC_57__cst_28__data__0__anchor__out = forkC_57_out1_data;
	assign cst_28_in1_valid = forkC_57__cst_28__valid__0__anchor__in;
	assign forkC_57__cst_28__valid__0__anchor__out = forkC_57_out1_valid;
	assign forkC_57_out1_ready = forkC_57__cst_28__ready__0__anchor__in;
	assign forkC_57__cst_28__ready__0__anchor__out = cst_28_in1_ready;
	assign branchC_59_in1_data = forkC_57__branchC_59__data__0__anchor__in;
	assign forkC_57__branchC_59__data__0__anchor__out = forkC_57_out2_data;
	assign branchC_59_in1_valid = forkC_57__branchC_59__valid__0__anchor__in;
	assign forkC_57__branchC_59__valid__0__anchor__out = forkC_57_out2_valid;
	assign forkC_57_out2_ready = forkC_57__branchC_59__ready__0__anchor__in;
	assign forkC_57__branchC_59__ready__0__anchor__out = branchC_59_in1_ready;
	assign branchC_59_clk = clk;
	assign branchC_59_rst = rst;
	assign Buffer_6_in1_data = branchC_59__Buffer_6__data__0__anchor__in;
	assign branchC_59__Buffer_6__data__0__anchor__out = branchC_59_out1_data;
	assign Buffer_6_in1_valid = branchC_59__Buffer_6__valid__0__anchor__in;
	assign branchC_59__Buffer_6__valid__0__anchor__out = branchC_59_out1_valid;
	assign branchC_59_out1_ready = branchC_59__Buffer_6__ready__0__anchor__in;
	assign branchC_59__Buffer_6__ready__0__anchor__out = Buffer_6_in1_ready;
	assign phiC_41_in1_data = branchC_59__phiC_41__data__0__anchor__in;
	assign branchC_59__phiC_41__data__0__anchor__out = branchC_59_out2_data;
	assign phiC_41_in1_valid = branchC_59__phiC_41__valid__0__anchor__in;
	assign branchC_59__phiC_41__valid__0__anchor__out = branchC_59_out2_valid;
	assign branchC_59_out2_ready = branchC_59__phiC_41__ready__0__anchor__in;
	assign branchC_59__phiC_41__ready__0__anchor__out = phiC_41_in1_ready;
	assign phiC_41_clk = clk;
	assign phiC_41_rst = rst;
	assign ret_0_in1_data = phiC_41__ret_0__data__0__anchor__in;
	assign phiC_41__ret_0__data__0__anchor__out = phiC_41_out1_data;
	assign ret_0_in1_valid = phiC_41__ret_0__valid__0__anchor__in;
	assign phiC_41__ret_0__valid__0__anchor__out = phiC_41_out1_valid;
	assign phiC_41_out1_ready = phiC_41__ret_0__ready__0__anchor__in;
	assign phiC_41__ret_0__ready__0__anchor__out = ret_0_in1_ready;
	assign sink_0_clk = clk;
	assign sink_0_rst = rst;
	assign sink_1_clk = clk;
	assign sink_1_rst = rst;
	assign sink_2_clk = clk;
	assign sink_2_rst = rst;
	assign sink_3_clk = clk;
	assign sink_3_rst = rst;
	assign sink_4_clk = clk;
	assign sink_4_rst = rst;
	assign sink_5_clk = clk;
	assign sink_5_rst = rst;
	assign sink_6_clk = clk;
	assign sink_6_rst = rst;
	assign sink_7_clk = clk;
	assign sink_7_rst = rst;
	assign sink_8_clk = clk;
	assign sink_8_rst = rst;
	assign sink_9_clk = clk;
	assign sink_9_rst = rst;
	assign sink_10_clk = clk;
	assign sink_10_rst = rst;
	assign sink_11_clk = clk;
	assign sink_11_rst = rst;
	assign sink_12_clk = clk;
	assign sink_12_rst = rst;
	assign sink_13_clk = clk;
	assign sink_13_rst = rst;
	assign sink_14_clk = clk;
	assign sink_14_rst = rst;
	assign sink_15_clk = clk;
	assign sink_15_rst = rst;
	assign sink_16_clk = clk;
	assign sink_16_rst = rst;
	assign sink_17_clk = clk;
	assign sink_17_rst = rst;
	assign sink_18_clk = clk;
	assign sink_18_rst = rst;
	assign sink_19_clk = clk;
	assign sink_19_rst = rst;
	assign sink_20_clk = clk;
	assign sink_20_rst = rst;
	assign sink_21_clk = clk;
	assign sink_21_rst = rst;
	assign sink_22_clk = clk;
	assign sink_22_rst = rst;
	assign sink_23_clk = clk;
	assign sink_23_rst = rst;
	assign sink_24_clk = clk;
	assign sink_24_rst = rst;
	assign sink_25_clk = clk;
	assign sink_25_rst = rst;
	assign sink_26_clk = clk;
	assign sink_26_rst = rst;
	assign sink_27_clk = clk;
	assign sink_27_rst = rst;
	assign sink_28_clk = clk;
	assign sink_28_rst = rst;
	assign sink_29_clk = clk;
	assign sink_29_rst = rst;
	assign sink_30_clk = clk;
	assign sink_30_rst = rst;
	assign sink_31_clk = clk;
	assign sink_31_rst = rst;
	assign sink_32_clk = clk;
	assign sink_32_rst = rst;
	assign sink_33_clk = clk;
	assign sink_33_rst = rst;
	assign sink_34_clk = clk;
	assign sink_34_rst = rst;
	assign sink_35_clk = clk;
	assign sink_35_rst = rst;
	assign sink_36_clk = clk;
	assign sink_36_rst = rst;
	assign sink_37_clk = clk;
	assign sink_37_rst = rst;
	assign sink_38_clk = clk;
	assign sink_38_rst = rst;
	assign source_0_clk = clk;
	assign source_0_rst = rst;
	assign cst_2_in1_data = source_0__cst_2__data__0__anchor__in;
	assign source_0__cst_2__data__0__anchor__out = source_0_out1_data;
	assign cst_2_in1_valid = source_0__cst_2__valid__0__anchor__in;
	assign source_0__cst_2__valid__0__anchor__out = source_0_out1_valid;
	assign source_0_out1_ready = source_0__cst_2__ready__0__anchor__in;
	assign source_0__cst_2__ready__0__anchor__out = cst_2_in1_ready;
	assign source_1_clk = clk;
	assign source_1_rst = rst;
	assign cst_3_in1_data = source_1__cst_3__data__0__anchor__in;
	assign source_1__cst_3__data__0__anchor__out = source_1_out1_data;
	assign cst_3_in1_valid = source_1__cst_3__valid__0__anchor__in;
	assign source_1__cst_3__valid__0__anchor__out = source_1_out1_valid;
	assign source_1_out1_ready = source_1__cst_3__ready__0__anchor__in;
	assign source_1__cst_3__ready__0__anchor__out = cst_3_in1_ready;
	assign source_2_clk = clk;
	assign source_2_rst = rst;
	assign cst_4_in1_data = source_2__cst_4__data__0__anchor__in;
	assign source_2__cst_4__data__0__anchor__out = source_2_out1_data;
	assign cst_4_in1_valid = source_2__cst_4__valid__0__anchor__in;
	assign source_2__cst_4__valid__0__anchor__out = source_2_out1_valid;
	assign source_2_out1_ready = source_2__cst_4__ready__0__anchor__in;
	assign source_2__cst_4__ready__0__anchor__out = cst_4_in1_ready;
	assign source_3_clk = clk;
	assign source_3_rst = rst;
	assign cst_5_in1_data = source_3__cst_5__data__0__anchor__in;
	assign source_3__cst_5__data__0__anchor__out = source_3_out1_data;
	assign cst_5_in1_valid = source_3__cst_5__valid__0__anchor__in;
	assign source_3__cst_5__valid__0__anchor__out = source_3_out1_valid;
	assign source_3_out1_ready = source_3__cst_5__ready__0__anchor__in;
	assign source_3__cst_5__ready__0__anchor__out = cst_5_in1_ready;
	assign source_4_clk = clk;
	assign source_4_rst = rst;
	assign cst_6_in1_data = source_4__cst_6__data__0__anchor__in;
	assign source_4__cst_6__data__0__anchor__out = source_4_out1_data;
	assign cst_6_in1_valid = source_4__cst_6__valid__0__anchor__in;
	assign source_4__cst_6__valid__0__anchor__out = source_4_out1_valid;
	assign source_4_out1_ready = source_4__cst_6__ready__0__anchor__in;
	assign source_4__cst_6__ready__0__anchor__out = cst_6_in1_ready;
	assign source_5_clk = clk;
	assign source_5_rst = rst;
	assign cst_7_in1_data = source_5__cst_7__data__0__anchor__in;
	assign source_5__cst_7__data__0__anchor__out = source_5_out1_data;
	assign cst_7_in1_valid = source_5__cst_7__valid__0__anchor__in;
	assign source_5__cst_7__valid__0__anchor__out = source_5_out1_valid;
	assign source_5_out1_ready = source_5__cst_7__ready__0__anchor__in;
	assign source_5__cst_7__ready__0__anchor__out = cst_7_in1_ready;
	assign source_6_clk = clk;
	assign source_6_rst = rst;
	assign cst_10_in1_data = source_6__cst_10__data__0__anchor__in;
	assign source_6__cst_10__data__0__anchor__out = source_6_out1_data;
	assign cst_10_in1_valid = source_6__cst_10__valid__0__anchor__in;
	assign source_6__cst_10__valid__0__anchor__out = source_6_out1_valid;
	assign source_6_out1_ready = source_6__cst_10__ready__0__anchor__in;
	assign source_6__cst_10__ready__0__anchor__out = cst_10_in1_ready;
	assign source_7_clk = clk;
	assign source_7_rst = rst;
	assign cst_11_in1_data = source_7__cst_11__data__0__anchor__in;
	assign source_7__cst_11__data__0__anchor__out = source_7_out1_data;
	assign cst_11_in1_valid = source_7__cst_11__valid__0__anchor__in;
	assign source_7__cst_11__valid__0__anchor__out = source_7_out1_valid;
	assign source_7_out1_ready = source_7__cst_11__ready__0__anchor__in;
	assign source_7__cst_11__ready__0__anchor__out = cst_11_in1_ready;
	assign source_8_clk = clk;
	assign source_8_rst = rst;
	assign cst_12_in1_data = source_8__cst_12__data__0__anchor__in;
	assign source_8__cst_12__data__0__anchor__out = source_8_out1_data;
	assign cst_12_in1_valid = source_8__cst_12__valid__0__anchor__in;
	assign source_8__cst_12__valid__0__anchor__out = source_8_out1_valid;
	assign source_8_out1_ready = source_8__cst_12__ready__0__anchor__in;
	assign source_8__cst_12__ready__0__anchor__out = cst_12_in1_ready;
	assign source_9_clk = clk;
	assign source_9_rst = rst;
	assign cst_13_in1_data = source_9__cst_13__data__0__anchor__in;
	assign source_9__cst_13__data__0__anchor__out = source_9_out1_data;
	assign cst_13_in1_valid = source_9__cst_13__valid__0__anchor__in;
	assign source_9__cst_13__valid__0__anchor__out = source_9_out1_valid;
	assign source_9_out1_ready = source_9__cst_13__ready__0__anchor__in;
	assign source_9__cst_13__ready__0__anchor__out = cst_13_in1_ready;
	assign source_10_clk = clk;
	assign source_10_rst = rst;
	assign cst_14_in1_data = source_10__cst_14__data__0__anchor__in;
	assign source_10__cst_14__data__0__anchor__out = source_10_out1_data;
	assign cst_14_in1_valid = source_10__cst_14__valid__0__anchor__in;
	assign source_10__cst_14__valid__0__anchor__out = source_10_out1_valid;
	assign source_10_out1_ready = source_10__cst_14__ready__0__anchor__in;
	assign source_10__cst_14__ready__0__anchor__out = cst_14_in1_ready;
	assign source_11_clk = clk;
	assign source_11_rst = rst;
	assign cst_16_in1_data = source_11__cst_16__data__0__anchor__in;
	assign source_11__cst_16__data__0__anchor__out = source_11_out1_data;
	assign cst_16_in1_valid = source_11__cst_16__valid__0__anchor__in;
	assign source_11__cst_16__valid__0__anchor__out = source_11_out1_valid;
	assign source_11_out1_ready = source_11__cst_16__ready__0__anchor__in;
	assign source_11__cst_16__ready__0__anchor__out = cst_16_in1_ready;
	assign source_12_clk = clk;
	assign source_12_rst = rst;
	assign cst_17_in1_data = source_12__cst_17__data__0__anchor__in;
	assign source_12__cst_17__data__0__anchor__out = source_12_out1_data;
	assign cst_17_in1_valid = source_12__cst_17__valid__0__anchor__in;
	assign source_12__cst_17__valid__0__anchor__out = source_12_out1_valid;
	assign source_12_out1_ready = source_12__cst_17__ready__0__anchor__in;
	assign source_12__cst_17__ready__0__anchor__out = cst_17_in1_ready;
	assign source_13_clk = clk;
	assign source_13_rst = rst;
	assign cst_20_in1_data = source_13__cst_20__data__0__anchor__in;
	assign source_13__cst_20__data__0__anchor__out = source_13_out1_data;
	assign cst_20_in1_valid = source_13__cst_20__valid__0__anchor__in;
	assign source_13__cst_20__valid__0__anchor__out = source_13_out1_valid;
	assign source_13_out1_ready = source_13__cst_20__ready__0__anchor__in;
	assign source_13__cst_20__ready__0__anchor__out = cst_20_in1_ready;
	assign source_14_clk = clk;
	assign source_14_rst = rst;
	assign cst_21_in1_data = source_14__cst_21__data__0__anchor__in;
	assign source_14__cst_21__data__0__anchor__out = source_14_out1_data;
	assign cst_21_in1_valid = source_14__cst_21__valid__0__anchor__in;
	assign source_14__cst_21__valid__0__anchor__out = source_14_out1_valid;
	assign source_14_out1_ready = source_14__cst_21__ready__0__anchor__in;
	assign source_14__cst_21__ready__0__anchor__out = cst_21_in1_ready;
	assign source_15_clk = clk;
	assign source_15_rst = rst;
	assign cst_22_in1_data = source_15__cst_22__data__0__anchor__in;
	assign source_15__cst_22__data__0__anchor__out = source_15_out1_data;
	assign cst_22_in1_valid = source_15__cst_22__valid__0__anchor__in;
	assign source_15__cst_22__valid__0__anchor__out = source_15_out1_valid;
	assign source_15_out1_ready = source_15__cst_22__ready__0__anchor__in;
	assign source_15__cst_22__ready__0__anchor__out = cst_22_in1_ready;
	assign source_16_clk = clk;
	assign source_16_rst = rst;
	assign cst_23_in1_data = source_16__cst_23__data__0__anchor__in;
	assign source_16__cst_23__data__0__anchor__out = source_16_out1_data;
	assign cst_23_in1_valid = source_16__cst_23__valid__0__anchor__in;
	assign source_16__cst_23__valid__0__anchor__out = source_16_out1_valid;
	assign source_16_out1_ready = source_16__cst_23__ready__0__anchor__in;
	assign source_16__cst_23__ready__0__anchor__out = cst_23_in1_ready;
	assign source_17_clk = clk;
	assign source_17_rst = rst;
	assign cst_24_in1_data = source_17__cst_24__data__0__anchor__in;
	assign source_17__cst_24__data__0__anchor__out = source_17_out1_data;
	assign cst_24_in1_valid = source_17__cst_24__valid__0__anchor__in;
	assign source_17__cst_24__valid__0__anchor__out = source_17_out1_valid;
	assign source_17_out1_ready = source_17__cst_24__ready__0__anchor__in;
	assign source_17__cst_24__ready__0__anchor__out = cst_24_in1_ready;
	assign fork_62_clk = clk;
	assign fork_62_rst = rst;
	assign phi_41_in1_data = fork_62__phi_41__data__0__anchor__in;
	assign fork_62__phi_41__data__0__anchor__out = fork_62_out1_data;
	assign phi_41_in1_valid = fork_62__phi_41__valid__0__anchor__in;
	assign fork_62__phi_41__valid__0__anchor__out = fork_62_out1_valid;
	assign fork_62_out1_ready = fork_62__phi_41__ready__0__anchor__in;
	assign fork_62__phi_41__ready__0__anchor__out = phi_41_in1_ready;
	assign phi_42_in1_data = fork_62__phi_42__data__0__anchor__in;
	assign fork_62__phi_42__data__0__anchor__out = fork_62_out2_data;
	assign phi_42_in1_valid = fork_62__phi_42__valid__0__anchor__in;
	assign fork_62__phi_42__valid__0__anchor__out = fork_62_out2_valid;
	assign fork_62_out2_ready = fork_62__phi_42__ready__0__anchor__in;
	assign fork_62__phi_42__ready__0__anchor__out = phi_42_in1_ready;
	assign fork_65_clk = clk;
	assign fork_65_rst = rst;
	assign phi_82_in1_data = fork_65__phi_82__data__0__anchor__in;
	assign fork_65__phi_82__data__0__anchor__out = fork_65_out1_data;
	assign phi_82_in1_valid = fork_65__phi_82__valid__0__anchor__in;
	assign fork_65__phi_82__valid__0__anchor__out = fork_65_out1_valid;
	assign fork_65_out1_ready = fork_65__phi_82__ready__0__anchor__in;
	assign fork_65__phi_82__ready__0__anchor__out = phi_82_in1_ready;
	assign phi_83_in1_data = fork_65__phi_83__data__0__anchor__in;
	assign fork_65__phi_83__data__0__anchor__out = fork_65_out2_data;
	assign phi_83_in1_valid = fork_65__phi_83__valid__0__anchor__in;
	assign fork_65__phi_83__valid__0__anchor__out = fork_65_out2_valid;
	assign fork_65_out2_ready = fork_65__phi_83__ready__0__anchor__in;
	assign fork_65__phi_83__ready__0__anchor__out = phi_83_in1_ready;
	assign Buffer_0_clk = clk;
	assign Buffer_0_rst = rst;
	assign phi_77_in3_data = Buffer_0__phi_77__data__0__anchor__in;
	assign Buffer_0__phi_77__data__0__anchor__out = Buffer_0_out1_data;
	assign phi_77_in3_valid = Buffer_0__phi_77__valid__0__anchor__in;
	assign Buffer_0__phi_77__valid__0__anchor__out = Buffer_0_out1_valid;
	assign Buffer_0_out1_ready = Buffer_0__phi_77__ready__0__anchor__in;
	assign Buffer_0__phi_77__ready__0__anchor__out = phi_77_in3_ready;
	assign Buffer_1_clk = clk;
	assign Buffer_1_rst = rst;
	assign phi_n0_in2_data = Buffer_1__phi_n0__data__0__anchor__in;
	assign Buffer_1__phi_n0__data__0__anchor__out = Buffer_1_out1_data;
	assign phi_n0_in2_valid = Buffer_1__phi_n0__valid__0__anchor__in;
	assign Buffer_1__phi_n0__valid__0__anchor__out = Buffer_1_out1_valid;
	assign Buffer_1_out1_ready = Buffer_1__phi_n0__ready__0__anchor__in;
	assign Buffer_1__phi_n0__ready__0__anchor__out = phi_n0_in2_ready;
	assign Buffer_2_clk = clk;
	assign Buffer_2_rst = rst;
	assign phiC_39_in2_data = Buffer_2__phiC_39__data__0__anchor__in;
	assign Buffer_2__phiC_39__data__0__anchor__out = Buffer_2_out1_data;
	assign phiC_39_in2_valid = Buffer_2__phiC_39__valid__0__anchor__in;
	assign Buffer_2__phiC_39__valid__0__anchor__out = Buffer_2_out1_valid;
	assign Buffer_2_out1_ready = Buffer_2__phiC_39__ready__0__anchor__in;
	assign Buffer_2__phiC_39__ready__0__anchor__out = phiC_39_in2_ready;
	assign Buffer_3_clk = clk;
	assign Buffer_3_rst = rst;
	assign phi_42_in3_data = Buffer_3__phi_42__data__0__anchor__in;
	assign Buffer_3__phi_42__data__0__anchor__out = Buffer_3_out1_data;
	assign phi_42_in3_valid = Buffer_3__phi_42__valid__0__anchor__in;
	assign Buffer_3__phi_42__valid__0__anchor__out = Buffer_3_out1_valid;
	assign Buffer_3_out1_ready = Buffer_3__phi_42__ready__0__anchor__in;
	assign Buffer_3__phi_42__ready__0__anchor__out = phi_42_in3_ready;
	assign Buffer_4_clk = clk;
	assign Buffer_4_rst = rst;
	assign phi_n6_in2_data = Buffer_4__phi_n6__data__0__anchor__in;
	assign Buffer_4__phi_n6__data__0__anchor__out = Buffer_4_out1_data;
	assign phi_n6_in2_valid = Buffer_4__phi_n6__valid__0__anchor__in;
	assign Buffer_4__phi_n6__valid__0__anchor__out = Buffer_4_out1_valid;
	assign Buffer_4_out1_ready = Buffer_4__phi_n6__ready__0__anchor__in;
	assign Buffer_4__phi_n6__ready__0__anchor__out = phi_n6_in2_ready;
	assign Buffer_5_clk = clk;
	assign Buffer_5_rst = rst;
	assign phi_n7_in2_data = Buffer_5__phi_n7__data__0__anchor__in;
	assign Buffer_5__phi_n7__data__0__anchor__out = Buffer_5_out1_data;
	assign phi_n7_in2_valid = Buffer_5__phi_n7__valid__0__anchor__in;
	assign Buffer_5__phi_n7__valid__0__anchor__out = Buffer_5_out1_valid;
	assign Buffer_5_out1_ready = Buffer_5__phi_n7__ready__0__anchor__in;
	assign Buffer_5__phi_n7__ready__0__anchor__out = phi_n7_in2_ready;
	assign Buffer_6_clk = clk;
	assign Buffer_6_rst = rst;
	assign phiC_38_in2_data = Buffer_6__phiC_38__data__0__anchor__in;
	assign Buffer_6__phiC_38__data__0__anchor__out = Buffer_6_out1_data;
	assign phiC_38_in2_valid = Buffer_6__phiC_38__valid__0__anchor__in;
	assign Buffer_6__phiC_38__valid__0__anchor__out = Buffer_6_out1_valid;
	assign Buffer_6_out1_ready = Buffer_6__phiC_38__ready__0__anchor__in;
	assign Buffer_6__phiC_38__ready__0__anchor__out = phiC_38_in2_ready;
	assign Buffer_7_clk = clk;
	assign Buffer_7_rst = rst;
	assign phiC_36_in2_data = Buffer_7__phiC_36__data__0__anchor__in;
	assign Buffer_7__phiC_36__data__0__anchor__out = Buffer_7_out1_data;
	assign phiC_36_in2_valid = Buffer_7__phiC_36__valid__0__anchor__in;
	assign Buffer_7__phiC_36__valid__0__anchor__out = Buffer_7_out1_valid;
	assign Buffer_7_out1_ready = Buffer_7__phiC_36__ready__0__anchor__in;
	assign Buffer_7__phiC_36__ready__0__anchor__out = phiC_36_in2_ready;
	assign Buffer_8_clk = clk;
	assign Buffer_8_rst = rst;
	assign phi_82_in3_data = Buffer_8__phi_82__data__0__anchor__in;
	assign Buffer_8__phi_82__data__0__anchor__out = Buffer_8_out1_data;
	assign phi_82_in3_valid = Buffer_8__phi_82__valid__0__anchor__in;
	assign Buffer_8__phi_82__valid__0__anchor__out = Buffer_8_out1_valid;
	assign Buffer_8_out1_ready = Buffer_8__phi_82__ready__0__anchor__in;
	assign Buffer_8__phi_82__ready__0__anchor__out = phi_82_in3_ready;
	assign Buffer_9_clk = clk;
	assign Buffer_9_rst = rst;
	assign phi_36_in3_data = Buffer_9__phi_36__data__0__anchor__in;
	assign Buffer_9__phi_36__data__0__anchor__out = Buffer_9_out1_data;
	assign phi_36_in3_valid = Buffer_9__phi_36__valid__0__anchor__in;
	assign Buffer_9__phi_36__valid__0__anchor__out = Buffer_9_out1_valid;
	assign Buffer_9_out1_ready = Buffer_9__phi_36__ready__0__anchor__in;
	assign Buffer_9__phi_36__ready__0__anchor__out = phi_36_in3_ready;
	assign Buffer_10_clk = clk;
	assign Buffer_10_rst = rst;
	assign phi_63_in3_data = Buffer_10__phi_63__data__0__anchor__in;
	assign Buffer_10__phi_63__data__0__anchor__out = Buffer_10_out1_data;
	assign phi_63_in3_valid = Buffer_10__phi_63__valid__0__anchor__in;
	assign Buffer_10__phi_63__valid__0__anchor__out = Buffer_10_out1_valid;
	assign Buffer_10_out1_ready = Buffer_10__phi_63__ready__0__anchor__in;
	assign Buffer_10__phi_63__ready__0__anchor__out = phi_63_in3_ready;
	assign Buffer_11_clk = clk;
	assign Buffer_11_rst = rst;
	assign phi_n22_in2_data = Buffer_11__phi_n22__data__0__anchor__in;
	assign Buffer_11__phi_n22__data__0__anchor__out = Buffer_11_out1_data;
	assign phi_n22_in2_valid = Buffer_11__phi_n22__valid__0__anchor__in;
	assign Buffer_11__phi_n22__valid__0__anchor__out = Buffer_11_out1_valid;
	assign Buffer_11_out1_ready = Buffer_11__phi_n22__ready__0__anchor__in;
	assign Buffer_11__phi_n22__ready__0__anchor__out = phi_n22_in2_ready;
	assign Buffer_12_clk = clk;
	assign Buffer_12_rst = rst;
	assign phi_41_in3_data = Buffer_12__phi_41__data__0__anchor__in;
	assign Buffer_12__phi_41__data__0__anchor__out = Buffer_12_out1_data;
	assign phi_41_in3_valid = Buffer_12__phi_41__valid__0__anchor__in;
	assign Buffer_12__phi_41__valid__0__anchor__out = Buffer_12_out1_valid;
	assign Buffer_12_out1_ready = Buffer_12__phi_41__ready__0__anchor__in;
	assign Buffer_12__phi_41__ready__0__anchor__out = phi_41_in3_ready;
	assign Buffer_13_clk = clk;
	assign Buffer_13_rst = rst;
	assign phi_n10_in2_data = Buffer_13__phi_n10__data__0__anchor__in;
	assign Buffer_13__phi_n10__data__0__anchor__out = Buffer_13_out1_data;
	assign phi_n10_in2_valid = Buffer_13__phi_n10__valid__0__anchor__in;
	assign Buffer_13__phi_n10__valid__0__anchor__out = Buffer_13_out1_valid;
	assign Buffer_13_out1_ready = Buffer_13__phi_n10__ready__0__anchor__in;
	assign Buffer_13__phi_n10__ready__0__anchor__out = phi_n10_in2_ready;
	assign Buffer_14_clk = clk;
	assign Buffer_14_rst = rst;
	assign phi_n5_in2_data = Buffer_14__phi_n5__data__0__anchor__in;
	assign Buffer_14__phi_n5__data__0__anchor__out = Buffer_14_out1_data;
	assign phi_n5_in2_valid = Buffer_14__phi_n5__valid__0__anchor__in;
	assign Buffer_14__phi_n5__valid__0__anchor__out = Buffer_14_out1_valid;
	assign Buffer_14_out1_ready = Buffer_14__phi_n5__ready__0__anchor__in;
	assign Buffer_14__phi_n5__ready__0__anchor__out = phi_n5_in2_ready;
	assign Buffer_15_clk = clk;
	assign Buffer_15_rst = rst;
	assign phi_n26_in2_data = Buffer_15__phi_n26__data__0__anchor__in;
	assign Buffer_15__phi_n26__data__0__anchor__out = Buffer_15_out1_data;
	assign phi_n26_in2_valid = Buffer_15__phi_n26__valid__0__anchor__in;
	assign Buffer_15__phi_n26__valid__0__anchor__out = Buffer_15_out1_valid;
	assign Buffer_15_out1_ready = Buffer_15__phi_n26__ready__0__anchor__in;
	assign Buffer_15__phi_n26__ready__0__anchor__out = phi_n26_in2_ready;
	assign Buffer_16_clk = clk;
	assign Buffer_16_rst = rst;
	assign phiC_28_in2_data = Buffer_16__phiC_28__data__0__anchor__in;
	assign Buffer_16__phiC_28__data__0__anchor__out = Buffer_16_out1_data;
	assign phiC_28_in2_valid = Buffer_16__phiC_28__valid__0__anchor__in;
	assign Buffer_16__phiC_28__valid__0__anchor__out = Buffer_16_out1_valid;
	assign Buffer_16_out1_ready = Buffer_16__phiC_28__ready__0__anchor__in;
	assign Buffer_16__phiC_28__ready__0__anchor__out = phiC_28_in2_ready;
	assign Buffer_17_clk = clk;
	assign Buffer_17_rst = rst;
	assign phi_n16_in2_data = Buffer_17__phi_n16__data__0__anchor__in;
	assign Buffer_17__phi_n16__data__0__anchor__out = Buffer_17_out1_data;
	assign phi_n16_in2_valid = Buffer_17__phi_n16__valid__0__anchor__in;
	assign Buffer_17__phi_n16__valid__0__anchor__out = Buffer_17_out1_valid;
	assign Buffer_17_out1_ready = Buffer_17__phi_n16__ready__0__anchor__in;
	assign Buffer_17__phi_n16__ready__0__anchor__out = phi_n16_in2_ready;
	assign Buffer_18_clk = clk;
	assign Buffer_18_rst = rst;
	assign phi_n18_in2_data = Buffer_18__phi_n18__data__0__anchor__in;
	assign Buffer_18__phi_n18__data__0__anchor__out = Buffer_18_out1_data;
	assign phi_n18_in2_valid = Buffer_18__phi_n18__valid__0__anchor__in;
	assign Buffer_18__phi_n18__valid__0__anchor__out = Buffer_18_out1_valid;
	assign Buffer_18_out1_ready = Buffer_18__phi_n18__ready__0__anchor__in;
	assign Buffer_18__phi_n18__ready__0__anchor__out = phi_n18_in2_ready;
	assign Buffer_19_clk = clk;
	assign Buffer_19_rst = rst;
	assign phi_n1_in2_data = Buffer_19__phi_n1__data__0__anchor__in;
	assign Buffer_19__phi_n1__data__0__anchor__out = Buffer_19_out1_data;
	assign phi_n1_in2_valid = Buffer_19__phi_n1__valid__0__anchor__in;
	assign Buffer_19__phi_n1__valid__0__anchor__out = Buffer_19_out1_valid;
	assign Buffer_19_out1_ready = Buffer_19__phi_n1__ready__0__anchor__in;
	assign Buffer_19__phi_n1__ready__0__anchor__out = phi_n1_in2_ready;
	assign Buffer_20_clk = clk;
	assign Buffer_20_rst = rst;
	assign phiC_29_in2_data = Buffer_20__phiC_29__data__0__anchor__in;
	assign Buffer_20__phiC_29__data__0__anchor__out = Buffer_20_out1_data;
	assign phiC_29_in2_valid = Buffer_20__phiC_29__valid__0__anchor__in;
	assign Buffer_20__phiC_29__valid__0__anchor__out = Buffer_20_out1_valid;
	assign Buffer_20_out1_ready = Buffer_20__phiC_29__ready__0__anchor__in;
	assign Buffer_20__phiC_29__ready__0__anchor__out = phiC_29_in2_ready;
	assign Buffer_21_clk = clk;
	assign Buffer_21_rst = rst;
	assign phiC_33_in2_data = Buffer_21__phiC_33__data__0__anchor__in;
	assign Buffer_21__phiC_33__data__0__anchor__out = Buffer_21_out1_data;
	assign phiC_33_in2_valid = Buffer_21__phiC_33__valid__0__anchor__in;
	assign Buffer_21__phiC_33__valid__0__anchor__out = Buffer_21_out1_valid;
	assign Buffer_21_out1_ready = Buffer_21__phiC_33__ready__0__anchor__in;
	assign Buffer_21__phiC_33__ready__0__anchor__out = phiC_33_in2_ready;
	assign Buffer_22_clk = clk;
	assign Buffer_22_rst = rst;
	assign phi_n17_in2_data = Buffer_22__phi_n17__data__0__anchor__in;
	assign Buffer_22__phi_n17__data__0__anchor__out = Buffer_22_out1_data;
	assign phi_n17_in2_valid = Buffer_22__phi_n17__valid__0__anchor__in;
	assign Buffer_22__phi_n17__valid__0__anchor__out = Buffer_22_out1_valid;
	assign Buffer_22_out1_ready = Buffer_22__phi_n17__ready__0__anchor__in;
	assign Buffer_22__phi_n17__ready__0__anchor__out = phi_n17_in2_ready;
	assign Buffer_23_clk = clk;
	assign Buffer_23_rst = rst;
	assign phi_n27_in2_data = Buffer_23__phi_n27__data__0__anchor__in;
	assign Buffer_23__phi_n27__data__0__anchor__out = Buffer_23_out1_data;
	assign phi_n27_in2_valid = Buffer_23__phi_n27__valid__0__anchor__in;
	assign Buffer_23__phi_n27__valid__0__anchor__out = Buffer_23_out1_valid;
	assign Buffer_23_out1_ready = Buffer_23__phi_n27__ready__0__anchor__in;
	assign Buffer_23__phi_n27__ready__0__anchor__out = phi_n27_in2_ready;
	assign Buffer_24_clk = clk;
	assign Buffer_24_rst = rst;
	assign phi_n11_in2_data = Buffer_24__phi_n11__data__0__anchor__in;
	assign Buffer_24__phi_n11__data__0__anchor__out = Buffer_24_out1_data;
	assign phi_n11_in2_valid = Buffer_24__phi_n11__valid__0__anchor__in;
	assign Buffer_24__phi_n11__valid__0__anchor__out = Buffer_24_out1_valid;
	assign Buffer_24_out1_ready = Buffer_24__phi_n11__ready__0__anchor__in;
	assign Buffer_24__phi_n11__ready__0__anchor__out = phi_n11_in2_ready;
	assign Buffer_25_clk = clk;
	assign Buffer_25_rst = rst;
	assign phi_3_in3_data = Buffer_25__phi_3__data__0__anchor__in;
	assign Buffer_25__phi_3__data__0__anchor__out = Buffer_25_out1_data;
	assign phi_3_in3_valid = Buffer_25__phi_3__valid__0__anchor__in;
	assign Buffer_25__phi_3__valid__0__anchor__out = Buffer_25_out1_valid;
	assign Buffer_25_out1_ready = Buffer_25__phi_3__ready__0__anchor__in;
	assign Buffer_25__phi_3__ready__0__anchor__out = phi_3_in3_ready;
	assign Buffer_26_clk = clk;
	assign Buffer_26_rst = rst;
	assign phi_1_in3_data = Buffer_26__phi_1__data__0__anchor__in;
	assign Buffer_26__phi_1__data__0__anchor__out = Buffer_26_out1_data;
	assign phi_1_in3_valid = Buffer_26__phi_1__valid__0__anchor__in;
	assign Buffer_26__phi_1__valid__0__anchor__out = Buffer_26_out1_valid;
	assign Buffer_26_out1_ready = Buffer_26__phi_1__ready__0__anchor__in;
	assign Buffer_26__phi_1__ready__0__anchor__out = phi_1_in3_ready;
	assign Buffer_27_clk = clk;
	assign Buffer_27_rst = rst;
	assign phiC_32_in2_data = Buffer_27__phiC_32__data__0__anchor__in;
	assign Buffer_27__phiC_32__data__0__anchor__out = Buffer_27_out1_data;
	assign phiC_32_in2_valid = Buffer_27__phiC_32__valid__0__anchor__in;
	assign Buffer_27__phiC_32__valid__0__anchor__out = Buffer_27_out1_valid;
	assign Buffer_27_out1_ready = Buffer_27__phiC_32__ready__0__anchor__in;
	assign Buffer_27__phiC_32__ready__0__anchor__out = phiC_32_in2_ready;
	assign Buffer_28_clk = clk;
	assign Buffer_28_rst = rst;
	assign phi_n20_in2_data = Buffer_28__phi_n20__data__0__anchor__in;
	assign Buffer_28__phi_n20__data__0__anchor__out = Buffer_28_out1_data;
	assign phi_n20_in2_valid = Buffer_28__phi_n20__valid__0__anchor__in;
	assign Buffer_28__phi_n20__valid__0__anchor__out = Buffer_28_out1_valid;
	assign Buffer_28_out1_ready = Buffer_28__phi_n20__ready__0__anchor__in;
	assign Buffer_28__phi_n20__ready__0__anchor__out = phi_n20_in2_ready;
	assign Buffer_29_clk = clk;
	assign Buffer_29_rst = rst;
	assign phi_83_in3_data = Buffer_29__phi_83__data__0__anchor__in;
	assign Buffer_29__phi_83__data__0__anchor__out = Buffer_29_out1_data;
	assign phi_83_in3_valid = Buffer_29__phi_83__valid__0__anchor__in;
	assign Buffer_29__phi_83__valid__0__anchor__out = Buffer_29_out1_valid;
	assign Buffer_29_out1_ready = Buffer_29__phi_83__ready__0__anchor__in;
	assign Buffer_29__phi_83__ready__0__anchor__out = phi_83_in3_ready;
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_32 (.clk(add_32_clk), .rst(add_32_rst), .data_in_bus({add_32_in2_data, add_32_in1_data}), .valid_in_bus({add_32_in2_valid, add_32_in1_valid}), .ready_in_bus({add_32_in2_ready, add_32_in1_ready}), .data_out_bus({add_32_out1_data}), .valid_out_bus({add_32_out1_valid}), .ready_out_bus({add_32_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_19 (.clk(sink_19_clk), .rst(sink_19_rst), .data_in_bus({sink_19_in1_data}), .valid_in_bus({sink_19_in1_valid}), .ready_in_bus({sink_19_in1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_26 (.clk(fork_26_clk), .rst(fork_26_rst), .data_in_bus({fork_26_in1_data}), .valid_in_bus({fork_26_in1_valid}), .ready_in_bus({fork_26_in1_ready}), .data_out_bus({fork_26_out2_data, fork_26_out1_data}), .valid_out_bus({fork_26_out2_valid, fork_26_out1_valid}), .ready_out_bus({fork_26_out2_ready, fork_26_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) OEHB_Buffer_3 (.clk(Buffer_3_clk), .rst(Buffer_3_rst), .data_in_bus({Buffer_3_in1_data}), .valid_in_bus({Buffer_3_in1_valid}), .ready_in_bus({Buffer_3_in1_ready}), .data_out_bus({Buffer_3_out1_data}), .valid_out_bus({Buffer_3_out1_valid}), .ready_out_bus({Buffer_3_out1_ready}));
shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(11), .DATA_OUT_SIZE(11)) shl_op_shl_43 (.clk(shl_43_clk), .rst(shl_43_rst), .data_in_bus({shl_43_in2_data, shl_43_in1_data}), .valid_in_bus({shl_43_in2_valid, shl_43_in1_valid}), .ready_in_bus({shl_43_in2_ready, shl_43_in1_ready}), .data_out_bus({shl_43_out1_data}), .valid_out_bus({shl_43_out1_valid}), .ready_out_bus({shl_43_out1_ready}));
icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_55 (.clk(icmp_55_clk), .rst(icmp_55_rst), .data_in_bus({icmp_55_in2_data, icmp_55_in1_data}), .valid_in_bus({icmp_55_in2_valid, icmp_55_in1_valid}), .ready_in_bus({icmp_55_in2_ready, icmp_55_in1_ready}), .data_out_bus({icmp_55_out1_data}), .valid_out_bus({icmp_55_out1_valid}), .ready_out_bus({icmp_55_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_11 (.clk(fork_11_clk), .rst(fork_11_rst), .data_in_bus({fork_11_in1_data}), .valid_in_bus({fork_11_in1_valid}), .ready_in_bus({fork_11_in1_ready}), .data_out_bus({fork_11_out3_data, fork_11_out2_data, fork_11_out1_data}), .valid_out_bus({fork_11_out3_valid, fork_11_out2_valid, fork_11_out1_valid}), .ready_out_bus({fork_11_out3_ready, fork_11_out2_ready, fork_11_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_28 (.clk(branch_28_clk), .rst(branch_28_rst), .data_in_bus({{5'b0, branch_28_in2_data}, branch_28_in1_data}), .valid_in_bus({branch_28_in2_valid, branch_28_in1_valid}), .ready_in_bus({branch_28_in2_ready, branch_28_in1_ready}), .data_out_bus({branch_28_out2_data, branch_28_out1_data}), .valid_out_bus({branch_28_out2_valid, branch_28_out1_valid}), .ready_out_bus({branch_28_out2_ready, branch_28_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) OEHB_Buffer_6 (.clk(Buffer_6_clk), .rst(Buffer_6_rst), .data_in_bus({Buffer_6_in1_data}), .valid_in_bus({Buffer_6_in1_valid}), .ready_in_bus({Buffer_6_in1_ready}), .data_out_bus({Buffer_6_out1_data}), .valid_out_bus({Buffer_6_out1_valid}), .ready_out_bus({Buffer_6_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_41 (.clk(branch_41_clk), .rst(branch_41_rst), .data_in_bus({{5'b0, branch_41_in2_data}, branch_41_in1_data}), .valid_in_bus({branch_41_in2_valid, branch_41_in1_valid}), .ready_in_bus({branch_41_in2_ready, branch_41_in1_ready}), .data_out_bus({branch_41_out2_data, branch_41_out1_data}), .valid_out_bus({branch_41_out2_valid, branch_41_out1_valid}), .ready_out_bus({branch_41_out2_ready, branch_41_out1_ready}));
cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_33 (.clk(phiC_33_clk), .rst(phiC_33_rst), .data_in_bus({phiC_33_in2_data, phiC_33_in1_data}), .valid_in_bus({phiC_33_in2_valid, phiC_33_in1_valid}), .ready_in_bus({phiC_33_in2_ready, phiC_33_in1_ready}), .data_out_bus({phiC_33_out2_data, phiC_33_out1_data}), .valid_out_bus({phiC_33_out2_valid, phiC_33_out1_valid}), .ready_out_bus({phiC_33_out2_ready, phiC_33_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_56 (.clk(branchC_56_clk), .rst(branchC_56_rst), .data_in_bus({{branchC_56_in2_data}, branchC_56_in1_data}), .valid_in_bus({branchC_56_in2_valid, branchC_56_in1_valid}), .ready_in_bus({branchC_56_in2_ready, branchC_56_in1_ready}), .data_out_bus({branchC_56_out2_data, branchC_56_out1_data}), .valid_out_bus({branchC_56_out2_valid, branchC_56_out1_valid}), .ready_out_bus({branchC_56_out2_ready, branchC_56_out1_ready}));
mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_36 (.clk(phi_36_clk), .rst(phi_36_rst), .data_in_bus({{5'b0, phi_36_in1_data}, phi_36_in3_data, phi_36_in2_data}), .valid_in_bus({phi_36_in1_valid, phi_36_in3_valid, phi_36_in2_valid}), .ready_in_bus({phi_36_in1_ready, phi_36_in3_ready, phi_36_in2_ready}), .data_out_bus({phi_36_out1_data}), .valid_out_bus({phi_36_out1_valid}), .ready_out_bus({phi_36_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_9 (.clk(fork_9_clk), .rst(fork_9_rst), .data_in_bus({fork_9_in1_data}), .valid_in_bus({fork_9_in1_valid}), .ready_in_bus({fork_9_in1_ready}), .data_out_bus({fork_9_out2_data, fork_9_out1_data}), .valid_out_bus({fork_9_out2_valid, fork_9_out1_valid}), .ready_out_bus({fork_9_out2_ready, fork_9_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_9 (.clk(sink_9_clk), .rst(sink_9_rst), .data_in_bus({sink_9_in1_data}), .valid_in_bus({sink_9_in1_valid}), .ready_in_bus({sink_9_in1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_39 (.clk(load_39_clk), .rst(load_39_rst), .data_in_bus({load_39_in1_data}), .address_in_bus({load_39_in2_data}), .valid_in_bus({load_39_in2_valid, load_39_in1_valid}), .ready_in_bus({load_39_in2_ready, load_39_in1_ready}), .data_out_bus({load_39_out1_data}), .address_out_bus({load_39_out2_data}), .valid_out_bus({load_39_out2_valid, load_39_out1_valid}), .ready_out_bus({load_39_out2_ready, load_39_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_48 (.clk(forkC_48_clk), .rst(forkC_48_rst), .data_in_bus({forkC_48_in1_data}), .valid_in_bus({forkC_48_in1_valid}), .ready_in_bus({forkC_48_in1_ready}), .data_out_bus({forkC_48_out3_data, forkC_48_out2_data, forkC_48_out1_data}), .valid_out_bus({forkC_48_out3_valid, forkC_48_out2_valid, forkC_48_out1_valid}), .ready_out_bus({forkC_48_out3_ready, forkC_48_out2_ready, forkC_48_out1_ready}));
start_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) start_node_beta (.clk(beta_clk), .rst(beta_rst), .data_in_bus({beta_in1_data}), .valid_in_bus({beta_in1_valid}), .ready_in_bus({beta_in1_ready}), .data_out_bus({beta_out1_data}), .valid_out_bus({beta_out1_valid}), .ready_out_bus({beta_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_34 (.clk(sink_34_clk), .rst(sink_34_rst), .data_in_bus({sink_34_in1_data}), .valid_in_bus({sink_34_in1_valid}), .ready_in_bus({sink_34_in1_ready}));
MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_y (.clk(MC_y_clk), .rst(MC_y_rst), .io_storeDataOut(y_dout0), .io_storeAddrOut(y_address0), .io_storeEnable(y_we0), .io_loadDataIn(y_din1), .io_loadAddrOut(y_address1), .io_loadEnable(y_ce1), .io_bbpValids({MC_y_in2_valid}), .io_bb_stCountArray({MC_y_in2_data}), .io_bbReadyToPrevs({MC_y_in2_ready}), .io_rdPortsPrev_ready({MC_y_in1_ready}), .io_rdPortsPrev_valid({MC_y_in1_valid}), .io_rdPortsPrev_bits({MC_y_in1_data}), .io_wrAddrPorts_ready({MC_y_in3_ready}), .io_wrAddrPorts_valid({MC_y_in3_valid}), .io_wrAddrPorts_bits({MC_y_in3_data}), .io_wrDataPorts_ready({MC_y_in4_ready}), .io_wrDataPorts_valid({MC_y_in4_valid}), .io_wrDataPorts_bits({MC_y_in4_data}), .io_rdPortsNext_ready({MC_y_out1_ready}), .io_rdPortsNext_valid({MC_y_out1_valid}), .io_rdPortsNext_bits({MC_y_out1_data}), .io_Empty_Valid({MC_y_out2_valid}), .io_Empty_Ready({MC_y_out2_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n14 (.clk(phi_n14_clk), .rst(phi_n14_rst), .data_in_bus({phi_n14_in1_data}), .valid_in_bus({phi_n14_in1_valid}), .ready_in_bus({phi_n14_in1_ready}), .data_out_bus({phi_n14_out1_data}), .valid_out_bus({phi_n14_out1_valid}), .ready_out_bus({phi_n14_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_80 (.clk(load_80_clk), .rst(load_80_rst), .data_in_bus({load_80_in1_data}), .address_in_bus({load_80_in2_data}), .valid_in_bus({load_80_in2_valid, load_80_in1_valid}), .ready_in_bus({load_80_in2_ready, load_80_in1_ready}), .data_out_bus({load_80_out1_data}), .address_out_bus({load_80_out2_data}), .valid_out_bus({load_80_out2_valid, load_80_out1_valid}), .ready_out_bus({load_80_out2_ready, load_80_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block1 (.clk(brCst_block1_clk), .rst(brCst_block1_rst), .data_in_bus({1'd1}), .valid_in_bus({brCst_block1_in1_valid}), .ready_in_bus({brCst_block1_in1_ready}), .data_out_bus({brCst_block1_out1_data}), .valid_out_bus({brCst_block1_out1_valid}), .ready_out_bus({brCst_block1_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_42 (.clk(fork_42_clk), .rst(fork_42_rst), .data_in_bus({fork_42_in1_data}), .valid_in_bus({fork_42_in1_valid}), .ready_in_bus({fork_42_in1_ready}), .data_out_bus({fork_42_out3_data, fork_42_out2_data, fork_42_out1_data}), .valid_out_bus({fork_42_out3_valid, fork_42_out2_valid, fork_42_out1_valid}), .ready_out_bus({fork_42_out3_ready, fork_42_out2_ready, fork_42_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n17 (.clk(phi_n17_clk), .rst(phi_n17_rst), .data_in_bus({phi_n17_in2_data, phi_n17_in1_data}), .valid_in_bus({phi_n17_in2_valid, phi_n17_in1_valid}), .ready_in_bus({phi_n17_in2_ready, phi_n17_in1_ready}), .data_out_bus({phi_n17_out1_data}), .valid_out_bus({phi_n17_out1_valid}), .ready_out_bus({phi_n17_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_2 (.clk(fork_2_clk), .rst(fork_2_rst), .data_in_bus({fork_2_in1_data}), .valid_in_bus({fork_2_in1_valid}), .ready_in_bus({fork_2_in1_ready}), .data_out_bus({fork_2_out2_data, fork_2_out1_data}), .valid_out_bus({fork_2_out2_valid, fork_2_out1_valid}), .ready_out_bus({fork_2_out2_ready, fork_2_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_36 (.clk(branch_36_clk), .rst(branch_36_rst), .data_in_bus({{31'b0, branch_36_in2_data}, branch_36_in1_data}), .valid_in_bus({branch_36_in2_valid, branch_36_in1_valid}), .ready_in_bus({branch_36_in2_ready, branch_36_in1_ready}), .data_out_bus({branch_36_out2_data, branch_36_out1_data}), .valid_out_bus({branch_36_out2_valid, branch_36_out1_valid}), .ready_out_bus({branch_36_out2_ready, branch_36_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_28 (.clk(sink_28_clk), .rst(sink_28_rst), .data_in_bus({sink_28_in1_data}), .valid_in_bus({sink_28_in1_valid}), .ready_in_bus({sink_28_in1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_1 (.clk(sink_1_clk), .rst(sink_1_rst), .data_in_bus({sink_1_in1_data}), .valid_in_bus({sink_1_in1_valid}), .ready_in_bus({sink_1_in1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(6), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_35 (.clk(fork_35_clk), .rst(fork_35_rst), .data_in_bus({fork_35_in1_data}), .valid_in_bus({fork_35_in1_valid}), .ready_in_bus({fork_35_in1_ready}), .data_out_bus({fork_35_out6_data, fork_35_out5_data, fork_35_out4_data, fork_35_out3_data, fork_35_out2_data, fork_35_out1_data}), .valid_out_bus({fork_35_out6_valid, fork_35_out5_valid, fork_35_out4_valid, fork_35_out3_valid, fork_35_out2_valid, fork_35_out1_valid}), .ready_out_bus({fork_35_out6_ready, fork_35_out5_ready, fork_35_out4_ready, fork_35_out3_ready, fork_35_out2_ready, fork_35_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_12 (.clk(sink_12_clk), .rst(sink_12_rst), .data_in_bus({sink_12_in1_data}), .valid_in_bus({sink_12_in1_valid}), .ready_in_bus({sink_12_in1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_13 (.clk(sink_13_clk), .rst(sink_13_rst), .data_in_bus({sink_13_in1_data}), .valid_in_bus({sink_13_in1_valid}), .ready_in_bus({sink_13_in1_ready}));
MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_z (.clk(MC_z_clk), .rst(MC_z_rst), .io_storeDataOut(z_dout0), .io_storeAddrOut(z_address0), .io_storeEnable(z_we0), .io_loadDataIn(z_din1), .io_loadAddrOut(z_address1), .io_loadEnable(z_ce1), .io_bbpValids({MC_z_in2_valid}), .io_bb_stCountArray({MC_z_in2_data}), .io_bbReadyToPrevs({MC_z_in2_ready}), .io_rdPortsPrev_ready({MC_z_in1_ready}), .io_rdPortsPrev_valid({MC_z_in1_valid}), .io_rdPortsPrev_bits({MC_z_in1_data}), .io_wrAddrPorts_ready({MC_z_in3_ready}), .io_wrAddrPorts_valid({MC_z_in3_valid}), .io_wrAddrPorts_bits({MC_z_in3_data}), .io_wrDataPorts_ready({MC_z_in4_ready}), .io_wrDataPorts_valid({MC_z_in4_valid}), .io_wrDataPorts_bits({MC_z_in4_data}), .io_rdPortsNext_ready({MC_z_out1_ready}), .io_rdPortsNext_valid({MC_z_out1_valid}), .io_rdPortsNext_bits({MC_z_out1_data}), .io_Empty_Valid({MC_z_out2_valid}), .io_Empty_Ready({MC_z_out2_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_7 (.clk(cst_7_clk), .rst(cst_7_rst), .data_in_bus({6'd32}), .valid_in_bus({cst_7_in1_valid}), .ready_in_bus({cst_7_in1_ready}), .data_out_bus({cst_7_out1_data}), .valid_out_bus({cst_7_out1_valid}), .ready_out_bus({cst_7_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block12 (.clk(brCst_block12_clk), .rst(brCst_block12_rst), .data_in_bus({1'd1}), .valid_in_bus({brCst_block12_in1_valid}), .ready_in_bus({brCst_block12_in1_ready}), .data_out_bus({brCst_block12_out1_data}), .valid_out_bus({brCst_block12_out1_valid}), .ready_out_bus({brCst_block12_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_18 (.clk(cst_18_clk), .rst(cst_18_rst), .data_in_bus({1'd0}), .valid_in_bus({cst_18_in1_valid}), .ready_in_bus({cst_18_in1_ready}), .data_out_bus({cst_18_out1_data}), .valid_out_bus({cst_18_out1_valid}), .ready_out_bus({cst_18_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_9 (.clk(cst_9_clk), .rst(cst_9_rst), .data_in_bus({1'd0}), .valid_in_bus({cst_9_in1_valid}), .ready_in_bus({cst_9_in1_ready}), .data_out_bus({cst_9_out1_data}), .valid_out_bus({cst_9_out1_valid}), .ready_out_bus({cst_9_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_32 (.clk(branch_32_clk), .rst(branch_32_rst), .data_in_bus({{5'b0, branch_32_in2_data}, branch_32_in1_data}), .valid_in_bus({branch_32_in2_valid, branch_32_in1_valid}), .ready_in_bus({branch_32_in2_ready, branch_32_in1_ready}), .data_out_bus({branch_32_out2_data, branch_32_out1_data}), .valid_out_bus({branch_32_out2_valid, branch_32_out1_valid}), .ready_out_bus({branch_32_out2_ready, branch_32_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_25 (.clk(sink_25_clk), .rst(sink_25_rst), .data_in_bus({sink_25_in1_data}), .valid_in_bus({sink_25_in1_valid}), .ready_in_bus({sink_25_in1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n22 (.clk(phi_n22_clk), .rst(phi_n22_rst), .data_in_bus({phi_n22_in2_data, phi_n22_in1_data}), .valid_in_bus({phi_n22_in2_valid, phi_n22_in1_valid}), .ready_in_bus({phi_n22_in2_ready, phi_n22_in1_ready}), .data_out_bus({phi_n22_out1_data}), .valid_out_bus({phi_n22_out1_valid}), .ready_out_bus({phi_n22_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) OEHB_Buffer_14 (.clk(Buffer_14_clk), .rst(Buffer_14_rst), .data_in_bus({Buffer_14_in1_data}), .valid_in_bus({Buffer_14_in1_valid}), .ready_in_bus({Buffer_14_in1_ready}), .data_out_bus({Buffer_14_out1_data}), .valid_out_bus({Buffer_14_out1_valid}), .ready_out_bus({Buffer_14_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_14 (.clk(cst_14_clk), .rst(cst_14_rst), .data_in_bus({6'd32}), .valid_in_bus({cst_14_in1_valid}), .ready_in_bus({cst_14_in1_ready}), .data_out_bus({cst_14_out1_data}), .valid_out_bus({cst_14_out1_valid}), .ready_out_bus({cst_14_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_6 (.clk(source_6_clk), .rst(source_6_rst), .data_out_bus({source_6_out1_data}), .valid_out_bus({source_6_out1_valid}), .ready_out_bus({source_6_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_4 (.clk(fork_4_clk), .rst(fork_4_rst), .data_in_bus({fork_4_in1_data}), .valid_in_bus({fork_4_in1_valid}), .ready_in_bus({fork_4_in1_ready}), .data_out_bus({fork_4_out3_data, fork_4_out2_data, fork_4_out1_data}), .valid_out_bus({fork_4_out3_valid, fork_4_out2_valid, fork_4_out1_valid}), .ready_out_bus({fork_4_out3_ready, fork_4_out2_ready, fork_4_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_38 (.clk(branch_38_clk), .rst(branch_38_rst), .data_in_bus({{31'b0, branch_38_in2_data}, branch_38_in1_data}), .valid_in_bus({branch_38_in2_valid, branch_38_in1_valid}), .ready_in_bus({branch_38_in2_ready, branch_38_in1_ready}), .data_out_bus({branch_38_out2_data, branch_38_out1_data}), .valid_out_bus({branch_38_out2_valid, branch_38_out1_valid}), .ready_out_bus({branch_38_out2_ready, branch_38_out1_ready}));
icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_101 (.clk(icmp_101_clk), .rst(icmp_101_rst), .data_in_bus({icmp_101_in2_data, icmp_101_in1_data}), .valid_in_bus({icmp_101_in2_valid, icmp_101_in1_valid}), .ready_in_bus({icmp_101_in2_ready, icmp_101_in1_ready}), .data_out_bus({icmp_101_out1_data}), .valid_out_bus({icmp_101_out1_valid}), .ready_out_bus({icmp_101_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_33 (.clk(sink_33_clk), .rst(sink_33_rst), .data_in_bus({sink_33_in1_data}), .valid_in_bus({sink_33_in1_valid}), .ready_in_bus({sink_33_in1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_43 (.clk(branch_43_clk), .rst(branch_43_rst), .data_in_bus({{31'b0, branch_43_in2_data}, branch_43_in1_data}), .valid_in_bus({branch_43_in2_valid, branch_43_in1_valid}), .ready_in_bus({branch_43_in2_ready, branch_43_in1_ready}), .data_out_bus({branch_43_out2_data, branch_43_out1_data}), .valid_out_bus({branch_43_out2_valid, branch_43_out1_valid}), .ready_out_bus({branch_43_out2_ready, branch_43_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n10 (.clk(phi_n10_clk), .rst(phi_n10_rst), .data_in_bus({phi_n10_in2_data, phi_n10_in1_data}), .valid_in_bus({phi_n10_in2_valid, phi_n10_in1_valid}), .ready_in_bus({phi_n10_in2_ready, phi_n10_in1_ready}), .data_out_bus({phi_n10_out1_data}), .valid_out_bus({phi_n10_out1_valid}), .ready_out_bus({phi_n10_out1_ready}));
mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(16), .DATA_OUT_SIZE(32)) mul_op_mul_52 (.clk(mul_52_clk), .rst(mul_52_rst), .data_in_bus({mul_52_in2_data, mul_52_in1_data}), .valid_in_bus({mul_52_in2_valid, mul_52_in1_valid}), .ready_in_bus({mul_52_in2_ready, mul_52_in1_ready}), .data_out_bus({mul_52_out1_data}), .valid_out_bus({mul_52_out1_valid}), .ready_out_bus({mul_52_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_20 (.clk(cst_20_clk), .rst(cst_20_rst), .data_in_bus({3'd5}), .valid_in_bus({cst_20_in1_valid}), .ready_in_bus({cst_20_in1_ready}), .data_out_bus({cst_20_out1_data}), .valid_out_bus({cst_20_out1_valid}), .ready_out_bus({cst_20_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_92 (.clk(load_92_clk), .rst(load_92_rst), .data_in_bus({load_92_in1_data}), .address_in_bus({load_92_in2_data}), .valid_in_bus({load_92_in2_valid, load_92_in1_valid}), .ready_in_bus({load_92_in2_ready, load_92_in1_ready}), .data_out_bus({load_92_out1_data}), .address_out_bus({load_92_out2_data}), .valid_out_bus({load_92_out2_valid, load_92_out1_valid}), .ready_out_bus({load_92_out2_ready, load_92_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_37 (.clk(sink_37_clk), .rst(sink_37_rst), .data_in_bus({sink_37_in1_data}), .valid_in_bus({sink_37_in1_valid}), .ready_in_bus({sink_37_in1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_17 (.clk(cst_17_clk), .rst(cst_17_rst), .data_in_bus({6'd32}), .valid_in_bus({cst_17_in1_valid}), .ready_in_bus({cst_17_in1_ready}), .data_out_bus({cst_17_out1_data}), .valid_out_bus({cst_17_out1_valid}), .ready_out_bus({cst_17_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) OEHB_Buffer_29 (.clk(Buffer_29_clk), .rst(Buffer_29_rst), .data_in_bus({Buffer_29_in1_data}), .valid_in_bus({Buffer_29_in1_valid}), .ready_in_bus({Buffer_29_in1_ready}), .data_out_bus({Buffer_29_out1_data}), .valid_out_bus({Buffer_29_out1_valid}), .ready_out_bus({Buffer_29_out1_ready}));
mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_3 (.clk(phi_3_clk), .rst(phi_3_rst), .data_in_bus({{5'b0, phi_3_in1_data}, phi_3_in3_data, phi_3_in2_data}), .valid_in_bus({phi_3_in1_valid, phi_3_in3_valid, phi_3_in2_valid}), .ready_in_bus({phi_3_in1_ready, phi_3_in3_ready, phi_3_in2_ready}), .data_out_bus({phi_3_out1_data}), .valid_out_bus({phi_3_out1_valid}), .ready_out_bus({phi_3_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_4 (.clk(Buffer_4_clk), .rst(Buffer_4_rst), .data_in_bus({Buffer_4_in1_data}), .valid_in_bus({Buffer_4_in1_valid}), .ready_in_bus({Buffer_4_in1_ready}), .data_out_bus({Buffer_4_out1_data}), .valid_out_bus({Buffer_4_out1_valid}), .ready_out_bus({Buffer_4_out1_ready}));
icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_60 (.clk(icmp_60_clk), .rst(icmp_60_rst), .data_in_bus({icmp_60_in2_data, icmp_60_in1_data}), .valid_in_bus({icmp_60_in2_valid, icmp_60_in1_valid}), .ready_in_bus({icmp_60_in2_ready, icmp_60_in1_ready}), .data_out_bus({icmp_60_out1_data}), .valid_out_bus({icmp_60_out1_valid}), .ready_out_bus({icmp_60_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_3 (.clk(sink_3_clk), .rst(sink_3_rst), .data_in_bus({sink_3_in1_data}), .valid_in_bus({sink_3_in1_valid}), .ready_in_bus({sink_3_in1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_5 (.clk(source_5_clk), .rst(source_5_rst), .data_out_bus({source_5_out1_data}), .valid_out_bus({source_5_out1_valid}), .ready_out_bus({source_5_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_18 (.clk(Buffer_18_clk), .rst(Buffer_18_rst), .data_in_bus({Buffer_18_in1_data}), .valid_in_bus({Buffer_18_in1_valid}), .ready_in_bus({Buffer_18_in1_ready}), .data_out_bus({Buffer_18_out1_data}), .valid_out_bus({Buffer_18_out1_valid}), .ready_out_bus({Buffer_18_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_49 (.clk(branchC_49_clk), .rst(branchC_49_rst), .data_in_bus({{branchC_49_in2_data}, branchC_49_in1_data}), .valid_in_bus({branchC_49_in2_valid, branchC_49_in1_valid}), .ready_in_bus({branchC_49_in2_ready, branchC_49_in1_ready}), .data_out_bus({branchC_49_out2_data, branchC_49_out1_data}), .valid_out_bus({branchC_49_out2_valid, branchC_49_out1_valid}), .ready_out_bus({branchC_49_out2_ready, branchC_49_out1_ready}));
mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(16), .DATA_OUT_SIZE(32)) mul_op_mul_93 (.clk(mul_93_clk), .rst(mul_93_rst), .data_in_bus({mul_93_in2_data, mul_93_in1_data}), .valid_in_bus({mul_93_in2_valid, mul_93_in1_valid}), .ready_in_bus({mul_93_in2_ready, mul_93_in1_ready}), .data_out_bus({mul_93_out1_data}), .valid_out_bus({mul_93_out1_valid}), .ready_out_bus({mul_93_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_11 (.clk(sink_11_clk), .rst(sink_11_rst), .data_in_bus({sink_11_in1_data}), .valid_in_bus({sink_11_in1_valid}), .ready_in_bus({sink_11_in1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_21 (.clk(sink_21_clk), .rst(sink_21_rst), .data_in_bus({sink_21_in1_data}), .valid_in_bus({sink_21_in1_valid}), .ready_in_bus({sink_21_in1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_22 (.clk(load_22_clk), .rst(load_22_rst), .data_in_bus({load_22_in1_data}), .address_in_bus({load_22_in2_data}), .valid_in_bus({load_22_in2_valid, load_22_in1_valid}), .ready_in_bus({load_22_in2_ready, load_22_in1_ready}), .data_out_bus({load_22_out1_data}), .address_out_bus({load_22_out2_data}), .valid_out_bus({load_22_out2_valid, load_22_out1_valid}), .ready_out_bus({load_22_out2_ready, load_22_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_28 (.clk(Buffer_28_clk), .rst(Buffer_28_rst), .data_in_bus({Buffer_28_in1_data}), .valid_in_bus({Buffer_28_in1_valid}), .ready_in_bus({Buffer_28_in1_ready}), .data_out_bus({Buffer_28_out1_data}), .valid_out_bus({Buffer_28_out1_valid}), .ready_out_bus({Buffer_28_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_45 (.clk(forkC_45_clk), .rst(forkC_45_rst), .data_in_bus({forkC_45_in1_data}), .valid_in_bus({forkC_45_in1_valid}), .ready_in_bus({forkC_45_in1_ready}), .data_out_bus({forkC_45_out3_data, forkC_45_out2_data, forkC_45_out1_data}), .valid_out_bus({forkC_45_out3_valid, forkC_45_out2_valid, forkC_45_out1_valid}), .ready_out_bus({forkC_45_out3_ready, forkC_45_out2_ready, forkC_45_out1_ready}));
end_node #(.INPUTS(1), .OUTPUTS(1), .MEMORY_INPUTS(9), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) end_node_end_0 (.clk(end_0_clk), .rst(end_0_rst), .data_in_bus({end_0_in10_data}), .valid_in_bus({end_0_in10_valid}), .ready_in_bus({end_0_in10_ready}), .e_valid_bus({end_0_in9_valid, end_0_in8_valid, end_0_in7_valid, end_0_in6_valid, end_0_in5_valid, end_0_in4_valid, end_0_in3_valid, end_0_in2_valid, end_0_in1_valid}), .e_ready_bus({end_0_in9_ready, end_0_in8_ready, end_0_in7_ready, end_0_in6_ready, end_0_in5_ready, end_0_in4_ready, end_0_in3_ready, end_0_in2_ready, end_0_in1_ready}), .data_out_bus({end_0_out1_data}), .valid_out_bus({end_0_out1_valid}), .ready_out_bus({end_0_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_59 (.clk(branchC_59_clk), .rst(branchC_59_rst), .data_in_bus({{branchC_59_in2_data}, branchC_59_in1_data}), .valid_in_bus({branchC_59_in2_valid, branchC_59_in1_valid}), .ready_in_bus({branchC_59_in2_ready, branchC_59_in1_ready}), .data_out_bus({branchC_59_out2_data, branchC_59_out1_data}), .valid_out_bus({branchC_59_out2_valid, branchC_59_out1_valid}), .ready_out_bus({branchC_59_out2_ready, branchC_59_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_10 (.clk(fork_10_clk), .rst(fork_10_rst), .data_in_bus({fork_10_in1_data}), .valid_in_bus({fork_10_in1_valid}), .ready_in_bus({fork_10_in1_ready}), .data_out_bus({fork_10_out2_data, fork_10_out1_data}), .valid_out_bus({fork_10_out2_valid, fork_10_out1_valid}), .ready_out_bus({fork_10_out2_ready, fork_10_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) OEHB_Buffer_9 (.clk(Buffer_9_clk), .rst(Buffer_9_rst), .data_in_bus({Buffer_9_in1_data}), .valid_in_bus({Buffer_9_in1_valid}), .ready_in_bus({Buffer_9_in1_ready}), .data_out_bus({Buffer_9_out1_data}), .valid_out_bus({Buffer_9_out1_valid}), .ready_out_bus({Buffer_9_out1_ready}));
cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_28 (.clk(phiC_28_clk), .rst(phiC_28_rst), .data_in_bus({phiC_28_in2_data, phiC_28_in1_data}), .valid_in_bus({phiC_28_in2_valid, phiC_28_in1_valid}), .ready_in_bus({phiC_28_in2_ready, phiC_28_in1_ready}), .data_out_bus({phiC_28_out2_data, phiC_28_out1_data}), .valid_out_bus({phiC_28_out2_valid, phiC_28_out1_valid}), .ready_out_bus({phiC_28_out2_ready, phiC_28_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_39 (.clk(fork_39_clk), .rst(fork_39_rst), .data_in_bus({fork_39_in1_data}), .valid_in_bus({fork_39_in1_valid}), .ready_in_bus({fork_39_in1_ready}), .data_out_bus({fork_39_out3_data, fork_39_out2_data, fork_39_out1_data}), .valid_out_bus({fork_39_out3_valid, fork_39_out2_valid, fork_39_out1_valid}), .ready_out_bus({fork_39_out3_ready, fork_39_out2_ready, fork_39_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_13 (.clk(Buffer_13_clk), .rst(Buffer_13_rst), .data_in_bus({Buffer_13_in1_data}), .valid_in_bus({Buffer_13_in1_valid}), .ready_in_bus({Buffer_13_in1_ready}), .data_out_bus({Buffer_13_out1_data}), .valid_out_bus({Buffer_13_out1_valid}), .ready_out_bus({Buffer_13_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_13 (.clk(fork_13_clk), .rst(fork_13_rst), .data_in_bus({fork_13_in1_data}), .valid_in_bus({fork_13_in1_valid}), .ready_in_bus({fork_13_in1_ready}), .data_out_bus({fork_13_out2_data, fork_13_out1_data}), .valid_out_bus({fork_13_out2_valid, fork_13_out1_valid}), .ready_out_bus({fork_13_out2_ready, fork_13_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_52 (.clk(forkC_52_clk), .rst(forkC_52_rst), .data_in_bus({forkC_52_in1_data}), .valid_in_bus({forkC_52_in1_valid}), .ready_in_bus({forkC_52_in1_ready}), .data_out_bus({forkC_52_out3_data, forkC_52_out2_data, forkC_52_out1_data}), .valid_out_bus({forkC_52_out3_valid, forkC_52_out2_valid, forkC_52_out1_valid}), .ready_out_bus({forkC_52_out3_ready, forkC_52_out2_ready, forkC_52_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) OEHB_Buffer_20 (.clk(Buffer_20_clk), .rst(Buffer_20_rst), .data_in_bus({Buffer_20_in1_data}), .valid_in_bus({Buffer_20_in1_valid}), .ready_in_bus({Buffer_20_in1_ready}), .data_out_bus({Buffer_20_out1_data}), .valid_out_bus({Buffer_20_out1_valid}), .ready_out_bus({Buffer_20_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_53 (.clk(branchC_53_clk), .rst(branchC_53_rst), .data_in_bus({{branchC_53_in2_data}, branchC_53_in1_data}), .valid_in_bus({branchC_53_in2_valid, branchC_53_in1_valid}), .ready_in_bus({branchC_53_in2_ready, branchC_53_in1_ready}), .data_out_bus({branchC_53_out2_data, branchC_53_out1_data}), .valid_out_bus({branchC_53_out2_valid, branchC_53_out1_valid}), .ready_out_bus({branchC_53_out2_ready, branchC_53_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_3 (.clk(source_3_clk), .rst(source_3_rst), .data_out_bus({source_3_out1_data}), .valid_out_bus({source_3_out1_valid}), .ready_out_bus({source_3_out1_ready}));
MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_w (.clk(MC_w_clk), .rst(MC_w_rst), .io_storeDataOut(w_dout0), .io_storeAddrOut(w_address0), .io_storeEnable(w_we0), .io_loadDataIn(w_din1), .io_loadAddrOut(w_address1), .io_loadEnable(w_ce1), .io_bbpValids({MC_w_in1_valid}), .io_bb_stCountArray({MC_w_in1_data}), .io_bbReadyToPrevs({MC_w_in1_ready}), .io_rdPortsPrev_ready({MC_w_in2_ready}), .io_rdPortsPrev_valid({MC_w_in2_valid}), .io_rdPortsPrev_bits({MC_w_in2_data}), .io_wrAddrPorts_ready({MC_w_in3_ready}), .io_wrAddrPorts_valid({MC_w_in3_valid}), .io_wrAddrPorts_bits({MC_w_in3_data}), .io_wrDataPorts_ready({MC_w_in4_ready}), .io_wrDataPorts_valid({MC_w_in4_valid}), .io_wrDataPorts_bits({MC_w_in4_data}), .io_rdPortsNext_ready({MC_w_out1_ready}), .io_rdPortsNext_valid({MC_w_out1_valid}), .io_rdPortsNext_bits({MC_w_out1_data}), .io_Empty_Valid({MC_w_out2_valid}), .io_Empty_Ready({MC_w_out2_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_24 (.clk(add_24_clk), .rst(add_24_rst), .data_in_bus({add_24_in2_data, add_24_in1_data}), .valid_in_bus({add_24_in2_valid, add_24_in1_valid}), .ready_in_bus({add_24_in2_ready, add_24_in1_ready}), .data_out_bus({add_24_out1_data}), .valid_out_bus({add_24_out1_valid}), .ready_out_bus({add_24_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_24 (.clk(Buffer_24_clk), .rst(Buffer_24_rst), .data_in_bus({Buffer_24_in1_data}), .valid_in_bus({Buffer_24_in1_valid}), .ready_in_bus({Buffer_24_in1_ready}), .data_out_bus({Buffer_24_out1_data}), .valid_out_bus({Buffer_24_out1_valid}), .ready_out_bus({Buffer_24_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_48 (.clk(branchC_48_clk), .rst(branchC_48_rst), .data_in_bus({{branchC_48_in2_data}, branchC_48_in1_data}), .valid_in_bus({branchC_48_in2_valid, branchC_48_in1_valid}), .ready_in_bus({branchC_48_in2_ready, branchC_48_in1_ready}), .data_out_bus({branchC_48_out2_data, branchC_48_out1_data}), .valid_out_bus({branchC_48_out2_valid, branchC_48_out1_valid}), .ready_out_bus({branchC_48_out2_ready, branchC_48_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_17 (.clk(fork_17_clk), .rst(fork_17_rst), .data_in_bus({fork_17_in1_data}), .valid_in_bus({fork_17_in1_valid}), .ready_in_bus({fork_17_in1_ready}), .data_out_bus({fork_17_out5_data, fork_17_out4_data, fork_17_out3_data, fork_17_out2_data, fork_17_out1_data}), .valid_out_bus({fork_17_out5_valid, fork_17_out4_valid, fork_17_out3_valid, fork_17_out2_valid, fork_17_out1_valid}), .ready_out_bus({fork_17_out5_ready, fork_17_out4_ready, fork_17_out3_ready, fork_17_out2_ready, fork_17_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n7 (.clk(phi_n7_clk), .rst(phi_n7_rst), .data_in_bus({phi_n7_in2_data, phi_n7_in1_data}), .valid_in_bus({phi_n7_in2_valid, phi_n7_in1_valid}), .ready_in_bus({phi_n7_in2_ready, phi_n7_in1_ready}), .data_out_bus({phi_n7_out1_data}), .valid_out_bus({phi_n7_out1_valid}), .ready_out_bus({phi_n7_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_4 (.clk(sink_4_clk), .rst(sink_4_rst), .data_in_bus({sink_4_in1_data}), .valid_in_bus({sink_4_in1_valid}), .ready_in_bus({sink_4_in1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) OEHB_Buffer_21 (.clk(Buffer_21_clk), .rst(Buffer_21_rst), .data_in_bus({Buffer_21_in1_data}), .valid_in_bus({Buffer_21_in1_valid}), .ready_in_bus({Buffer_21_in1_ready}), .data_out_bus({Buffer_21_out1_data}), .valid_out_bus({Buffer_21_out1_valid}), .ready_out_bus({Buffer_21_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_65 (.clk(fork_65_clk), .rst(fork_65_rst), .data_in_bus({fork_65_in1_data}), .valid_in_bus({fork_65_in1_valid}), .ready_in_bus({fork_65_in1_ready}), .data_out_bus({fork_65_out2_data, fork_65_out1_data}), .valid_out_bus({fork_65_out2_valid, fork_65_out1_valid}), .ready_out_bus({fork_65_out2_ready, fork_65_out1_ready}));
mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(16), .DATA_OUT_SIZE(32)) mul_op_mul_23 (.clk(mul_23_clk), .rst(mul_23_rst), .data_in_bus({mul_23_in2_data, mul_23_in1_data}), .valid_in_bus({mul_23_in2_valid, mul_23_in1_valid}), .ready_in_bus({mul_23_in2_ready, mul_23_in1_ready}), .data_out_bus({mul_23_out1_data}), .valid_out_bus({mul_23_out1_valid}), .ready_out_bus({mul_23_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_30 (.clk(fork_30_clk), .rst(fork_30_rst), .data_in_bus({fork_30_in1_data}), .valid_in_bus({fork_30_in1_valid}), .ready_in_bus({fork_30_in1_ready}), .data_out_bus({fork_30_out5_data, fork_30_out4_data, fork_30_out3_data, fork_30_out2_data, fork_30_out1_data}), .valid_out_bus({fork_30_out5_valid, fork_30_out4_valid, fork_30_out3_valid, fork_30_out2_valid, fork_30_out1_valid}), .ready_out_bus({fork_30_out5_ready, fork_30_out4_ready, fork_30_out3_ready, fork_30_out2_ready, fork_30_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_16 (.clk(source_16_clk), .rst(source_16_rst), .data_out_bus({source_16_out1_data}), .valid_out_bus({source_16_out1_valid}), .ready_out_bus({source_16_out1_ready}));
start_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) start_node_start_0 (.clk(start_0_clk), .rst(start_0_rst), .data_in_bus({start_0_in1_data}), .valid_in_bus({start_0_in1_valid}), .ready_in_bus({start_0_in1_ready}), .data_out_bus({start_0_out1_data}), .valid_out_bus({start_0_out1_valid}), .ready_out_bus({start_0_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) OEHB_Buffer_17 (.clk(Buffer_17_clk), .rst(Buffer_17_rst), .data_in_bus({Buffer_17_in1_data}), .valid_in_bus({Buffer_17_in1_valid}), .ready_in_bus({Buffer_17_in1_ready}), .data_out_bus({Buffer_17_out1_data}), .valid_out_bus({Buffer_17_out1_valid}), .ready_out_bus({Buffer_17_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_30 (.clk(branch_30_clk), .rst(branch_30_rst), .data_in_bus({{branch_30_in2_data}, branch_30_in1_data}), .valid_in_bus({branch_30_in2_valid, branch_30_in1_valid}), .ready_in_bus({branch_30_in2_ready, branch_30_in1_ready}), .data_out_bus({branch_30_out2_data, branch_30_out1_data}), .valid_out_bus({branch_30_out2_valid, branch_30_out1_valid}), .ready_out_bus({branch_30_out2_ready, branch_30_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_7 (.clk(branch_7_clk), .rst(branch_7_rst), .data_in_bus({{5'b0, branch_7_in2_data}, branch_7_in1_data}), .valid_in_bus({branch_7_in2_valid, branch_7_in1_valid}), .ready_in_bus({branch_7_in2_ready, branch_7_in1_ready}), .data_out_bus({branch_7_out2_data, branch_7_out1_data}), .valid_out_bus({branch_7_out2_valid, branch_7_out1_valid}), .ready_out_bus({branch_7_out2_ready, branch_7_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(12), .DATA_SIZE(32)) mc_load_op_load_8 (.clk(load_8_clk), .rst(load_8_rst), .data_in_bus({load_8_in1_data}), .address_in_bus({load_8_in2_data}), .valid_in_bus({load_8_in2_valid, load_8_in1_valid}), .ready_in_bus({load_8_in2_ready, load_8_in1_ready}), .data_out_bus({load_8_out1_data}), .address_out_bus({load_8_out2_data}), .valid_out_bus({load_8_out2_valid, load_8_out1_valid}), .ready_out_bus({load_8_out2_ready, load_8_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_22 (.clk(Buffer_22_clk), .rst(Buffer_22_rst), .data_in_bus({Buffer_22_in1_data}), .valid_in_bus({Buffer_22_in1_valid}), .ready_in_bus({Buffer_22_in1_ready}), .data_out_bus({Buffer_22_out1_data}), .valid_out_bus({Buffer_22_out1_valid}), .ready_out_bus({Buffer_22_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_20 (.clk(branch_20_clk), .rst(branch_20_rst), .data_in_bus({{31'b0, branch_20_in2_data}, branch_20_in1_data}), .valid_in_bus({branch_20_in2_valid, branch_20_in1_valid}), .ready_in_bus({branch_20_in2_ready, branch_20_in1_ready}), .data_out_bus({branch_20_out2_data, branch_20_out1_data}), .valid_out_bus({branch_20_out2_valid, branch_20_out1_valid}), .ready_out_bus({branch_20_out2_ready, branch_20_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_35 (.clk(branch_35_clk), .rst(branch_35_rst), .data_in_bus({{31'b0, branch_35_in2_data}, branch_35_in1_data}), .valid_in_bus({branch_35_in2_valid, branch_35_in1_valid}), .ready_in_bus({branch_35_in2_ready, branch_35_in1_ready}), .data_out_bus({branch_35_out2_data, branch_35_out1_data}), .valid_out_bus({branch_35_out2_valid, branch_35_out1_valid}), .ready_out_bus({branch_35_out2_ready, branch_35_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_38 (.clk(fork_38_clk), .rst(fork_38_rst), .data_in_bus({fork_38_in1_data}), .valid_in_bus({fork_38_in1_valid}), .ready_in_bus({fork_38_in1_ready}), .data_out_bus({fork_38_out3_data, fork_38_out2_data, fork_38_out1_data}), .valid_out_bus({fork_38_out3_valid, fork_38_out2_valid, fork_38_out1_valid}), .ready_out_bus({fork_38_out3_ready, fork_38_out2_ready, fork_38_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_6 (.clk(branch_6_clk), .rst(branch_6_rst), .data_in_bus({{31'b0, branch_6_in2_data}, branch_6_in1_data}), .valid_in_bus({branch_6_in2_valid, branch_6_in1_valid}), .ready_in_bus({branch_6_in2_ready, branch_6_in1_ready}), .data_out_bus({branch_6_out2_data, branch_6_out1_data}), .valid_out_bus({branch_6_out2_valid, branch_6_out1_valid}), .ready_out_bus({branch_6_out2_ready, branch_6_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_30 (.clk(Buffer_30_clk), .rst(Buffer_30_rst), .data_in_bus({Buffer_30_in1_data}), .valid_in_bus({Buffer_30_in1_valid}), .ready_in_bus({Buffer_30_in1_ready}), .data_out_bus({Buffer_30_out1_data}), .valid_out_bus({Buffer_30_out1_valid}), .ready_out_bus({Buffer_30_out1_ready}));
mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_42 (.clk(phi_42_clk), .rst(phi_42_rst), .data_in_bus({{5'b0, phi_42_in1_data}, phi_42_in3_data, phi_42_in2_data}), .valid_in_bus({phi_42_in1_valid, phi_42_in3_valid, phi_42_in2_valid}), .ready_in_bus({phi_42_in1_ready, phi_42_in3_ready, phi_42_in2_ready}), .data_out_bus({phi_42_out1_data}), .valid_out_bus({phi_42_out1_valid}), .ready_out_bus({phi_42_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_28 (.clk(fork_28_clk), .rst(fork_28_rst), .data_in_bus({fork_28_in1_data}), .valid_in_bus({fork_28_in1_valid}), .ready_in_bus({fork_28_in1_ready}), .data_out_bus({fork_28_out2_data, fork_28_out1_data}), .valid_out_bus({fork_28_out2_valid, fork_28_out1_valid}), .ready_out_bus({fork_28_out2_ready, fork_28_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n15 (.clk(phi_n15_clk), .rst(phi_n15_rst), .data_in_bus({phi_n15_in1_data}), .valid_in_bus({phi_n15_in1_valid}), .ready_in_bus({phi_n15_in1_ready}), .data_out_bus({phi_n15_out1_data}), .valid_out_bus({phi_n15_out1_valid}), .ready_out_bus({phi_n15_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_7 (.clk(source_7_clk), .rst(source_7_rst), .data_out_bus({source_7_out1_data}), .valid_out_bus({source_7_out1_valid}), .ready_out_bus({source_7_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_21 (.clk(branch_21_clk), .rst(branch_21_rst), .data_in_bus({{5'b0, branch_21_in2_data}, branch_21_in1_data}), .valid_in_bus({branch_21_in2_valid, branch_21_in1_valid}), .ready_in_bus({branch_21_in2_ready, branch_21_in1_ready}), .data_out_bus({branch_21_out2_data, branch_21_out1_data}), .valid_out_bus({branch_21_out2_valid, branch_21_out1_valid}), .ready_out_bus({branch_21_out2_ready, branch_21_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n4 (.clk(phi_n4_clk), .rst(phi_n4_rst), .data_in_bus({phi_n4_in1_data}), .valid_in_bus({phi_n4_in1_valid}), .ready_in_bus({phi_n4_in1_ready}), .data_out_bus({phi_n4_out1_data}), .valid_out_bus({phi_n4_out1_valid}), .ready_out_bus({phi_n4_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_53 (.clk(add_53_clk), .rst(add_53_rst), .data_in_bus({add_53_in2_data, add_53_in1_data}), .valid_in_bus({add_53_in2_valid, add_53_in1_valid}), .ready_in_bus({add_53_in2_ready, add_53_in1_ready}), .data_out_bus({add_53_out1_data}), .valid_out_bus({add_53_out1_valid}), .ready_out_bus({add_53_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_10 (.clk(cst_10_clk), .rst(cst_10_rst), .data_in_bus({3'd5}), .valid_in_bus({cst_10_in1_valid}), .ready_in_bus({cst_10_in1_ready}), .data_out_bus({cst_10_out1_data}), .valid_out_bus({cst_10_out1_valid}), .ready_out_bus({cst_10_out1_ready}));
icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_96 (.clk(icmp_96_clk), .rst(icmp_96_rst), .data_in_bus({icmp_96_in2_data, icmp_96_in1_data}), .valid_in_bus({icmp_96_in2_valid, icmp_96_in1_valid}), .ready_in_bus({icmp_96_in2_ready, icmp_96_in1_ready}), .data_out_bus({icmp_96_out1_data}), .valid_out_bus({icmp_96_out1_valid}), .ready_out_bus({icmp_96_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_7 (.clk(fork_7_clk), .rst(fork_7_rst), .data_in_bus({fork_7_in1_data}), .valid_in_bus({fork_7_in1_valid}), .ready_in_bus({fork_7_in1_ready}), .data_out_bus({fork_7_out2_data, fork_7_out1_data}), .valid_out_bus({fork_7_out2_valid, fork_7_out1_valid}), .ready_out_bus({fork_7_out2_ready, fork_7_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_55 (.clk(forkC_55_clk), .rst(forkC_55_rst), .data_in_bus({forkC_55_in1_data}), .valid_in_bus({forkC_55_in1_valid}), .ready_in_bus({forkC_55_in1_ready}), .data_out_bus({forkC_55_out3_data, forkC_55_out2_data, forkC_55_out1_data}), .valid_out_bus({forkC_55_out3_valid, forkC_55_out2_valid, forkC_55_out1_valid}), .ready_out_bus({forkC_55_out3_ready, forkC_55_out2_ready, forkC_55_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_33 (.clk(branch_33_clk), .rst(branch_33_rst), .data_in_bus({{31'b0, branch_33_in2_data}, branch_33_in1_data}), .valid_in_bus({branch_33_in2_valid, branch_33_in1_valid}), .ready_in_bus({branch_33_in2_ready, branch_33_in1_ready}), .data_out_bus({branch_33_out2_data, branch_33_out1_data}), .valid_out_bus({branch_33_out2_valid, branch_33_out1_valid}), .ready_out_bus({branch_33_out2_ready, branch_33_out1_ready}));
cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_29 (.clk(phiC_29_clk), .rst(phiC_29_rst), .data_in_bus({phiC_29_in2_data, phiC_29_in1_data}), .valid_in_bus({phiC_29_in2_valid, phiC_29_in1_valid}), .ready_in_bus({phiC_29_in2_ready, phiC_29_in1_ready}), .data_out_bus({phiC_29_out2_data, phiC_29_out1_data}), .valid_out_bus({phiC_29_out2_valid, phiC_29_out1_valid}), .ready_out_bus({phiC_29_out2_ready, phiC_29_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_46 (.clk(forkC_46_clk), .rst(forkC_46_rst), .data_in_bus({forkC_46_in1_data}), .valid_in_bus({forkC_46_in1_valid}), .ready_in_bus({forkC_46_in1_ready}), .data_out_bus({forkC_46_out2_data, forkC_46_out1_data}), .valid_out_bus({forkC_46_out2_valid, forkC_46_out1_valid}), .ready_out_bus({forkC_46_out2_ready, forkC_46_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_24 (.clk(branch_24_clk), .rst(branch_24_rst), .data_in_bus({{5'b0, branch_24_in2_data}, branch_24_in1_data}), .valid_in_bus({branch_24_in2_valid, branch_24_in1_valid}), .ready_in_bus({branch_24_in2_ready, branch_24_in1_ready}), .data_out_bus({branch_24_out2_data, branch_24_out1_data}), .valid_out_bus({branch_24_out2_valid, branch_24_out1_valid}), .ready_out_bus({branch_24_out2_ready, branch_24_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_22 (.clk(cst_22_clk), .rst(cst_22_rst), .data_in_bus({6'd32}), .valid_in_bus({cst_22_in1_valid}), .ready_in_bus({cst_22_in1_ready}), .data_out_bus({cst_22_out1_data}), .valid_out_bus({cst_22_out1_valid}), .ready_out_bus({cst_22_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_35 (.clk(sink_35_clk), .rst(sink_35_rst), .data_in_bus({sink_35_in1_data}), .valid_in_bus({sink_35_in1_valid}), .ready_in_bus({sink_35_in1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n11 (.clk(phi_n11_clk), .rst(phi_n11_rst), .data_in_bus({phi_n11_in2_data, phi_n11_in1_data}), .valid_in_bus({phi_n11_in2_valid, phi_n11_in1_valid}), .ready_in_bus({phi_n11_in2_ready, phi_n11_in1_ready}), .data_out_bus({phi_n11_out1_data}), .valid_out_bus({phi_n11_out1_valid}), .ready_out_bus({phi_n11_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_38 (.clk(sink_38_clk), .rst(sink_38_rst), .data_in_bus({sink_38_in1_data}), .valid_in_bus({sink_38_in1_valid}), .ready_in_bus({sink_38_in1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_40 (.clk(fork_40_clk), .rst(fork_40_rst), .data_in_bus({fork_40_in1_data}), .valid_in_bus({fork_40_in1_valid}), .ready_in_bus({fork_40_in1_ready}), .data_out_bus({fork_40_out5_data, fork_40_out4_data, fork_40_out3_data, fork_40_out2_data, fork_40_out1_data}), .valid_out_bus({fork_40_out5_valid, fork_40_out4_valid, fork_40_out3_valid, fork_40_out2_valid, fork_40_out1_valid}), .ready_out_bus({fork_40_out5_ready, fork_40_out4_ready, fork_40_out3_ready, fork_40_out2_ready, fork_40_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_62 (.clk(fork_62_clk), .rst(fork_62_rst), .data_in_bus({fork_62_in1_data}), .valid_in_bus({fork_62_in1_valid}), .ready_in_bus({fork_62_in1_ready}), .data_out_bus({fork_62_out2_data, fork_62_out1_data}), .valid_out_bus({fork_62_out2_valid, fork_62_out1_valid}), .ready_out_bus({fork_62_out2_ready, fork_62_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_57 (.clk(forkC_57_clk), .rst(forkC_57_rst), .data_in_bus({forkC_57_in1_data}), .valid_in_bus({forkC_57_in1_valid}), .ready_in_bus({forkC_57_in1_ready}), .data_out_bus({forkC_57_out2_data, forkC_57_out1_data}), .valid_out_bus({forkC_57_out2_valid, forkC_57_out1_valid}), .ready_out_bus({forkC_57_out2_ready, forkC_57_out1_ready}));
mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(16), .DATA_OUT_SIZE(32)) mul_op_mul_15 (.clk(mul_15_clk), .rst(mul_15_rst), .data_in_bus({mul_15_in2_data, mul_15_in1_data}), .valid_in_bus({mul_15_in2_valid, mul_15_in1_valid}), .ready_in_bus({mul_15_in2_ready, mul_15_in1_ready}), .data_out_bus({mul_15_out1_data}), .valid_out_bus({mul_15_out1_valid}), .ready_out_bus({mul_15_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_37 (.clk(fork_37_clk), .rst(fork_37_rst), .data_in_bus({fork_37_in1_data}), .valid_in_bus({fork_37_in1_valid}), .ready_in_bus({fork_37_in1_ready}), .data_out_bus({fork_37_out3_data, fork_37_out2_data, fork_37_out1_data}), .valid_out_bus({fork_37_out3_valid, fork_37_out2_valid, fork_37_out1_valid}), .ready_out_bus({fork_37_out3_ready, fork_37_out2_ready, fork_37_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(12), .DATA_OUT_SIZE(12)) add_op_add_44 (.clk(add_44_clk), .rst(add_44_rst), .data_in_bus({add_44_in2_data, add_44_in1_data}), .valid_in_bus({add_44_in2_valid, add_44_in1_valid}), .ready_in_bus({add_44_in2_ready, add_44_in1_ready}), .data_out_bus({add_44_out1_data}), .valid_out_bus({add_44_out1_valid}), .ready_out_bus({add_44_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_8 (.clk(fork_8_clk), .rst(fork_8_rst), .data_in_bus({fork_8_in1_data}), .valid_in_bus({fork_8_in1_valid}), .ready_in_bus({fork_8_in1_ready}), .data_out_bus({fork_8_out4_data, fork_8_out3_data, fork_8_out2_data, fork_8_out1_data}), .valid_out_bus({fork_8_out4_valid, fork_8_out3_valid, fork_8_out2_valid, fork_8_out1_valid}), .ready_out_bus({fork_8_out4_ready, fork_8_out3_ready, fork_8_out2_ready, fork_8_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n0 (.clk(phi_n0_clk), .rst(phi_n0_rst), .data_in_bus({phi_n0_in2_data, phi_n0_in1_data}), .valid_in_bus({phi_n0_in2_valid, phi_n0_in1_valid}), .ready_in_bus({phi_n0_in2_ready, phi_n0_in1_ready}), .data_out_bus({phi_n0_out1_data}), .valid_out_bus({phi_n0_out1_valid}), .ready_out_bus({phi_n0_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_4 (.clk(cst_4_clk), .rst(cst_4_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_4_in1_valid}), .ready_in_bus({cst_4_in1_ready}), .data_out_bus({cst_4_out1_data}), .valid_out_bus({cst_4_out1_valid}), .ready_out_bus({cst_4_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_25 (.clk(cst_25_clk), .rst(cst_25_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_25_in1_valid}), .ready_in_bus({cst_25_in1_ready}), .data_out_bus({cst_25_out1_data}), .valid_out_bus({cst_25_out1_valid}), .ready_out_bus({cst_25_out1_ready}));
icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_30 (.clk(icmp_30_clk), .rst(icmp_30_rst), .data_in_bus({icmp_30_in2_data, icmp_30_in1_data}), .valid_in_bus({icmp_30_in2_valid, icmp_30_in1_valid}), .ready_in_bus({icmp_30_in2_ready, icmp_30_in1_ready}), .data_out_bus({icmp_30_out1_data}), .valid_out_bus({icmp_30_out1_valid}), .ready_out_bus({icmp_30_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) OEHB_Buffer_15 (.clk(Buffer_15_clk), .rst(Buffer_15_rst), .data_in_bus({Buffer_15_in1_data}), .valid_in_bus({Buffer_15_in1_valid}), .ready_in_bus({Buffer_15_in1_ready}), .data_out_bus({Buffer_15_out1_data}), .valid_out_bus({Buffer_15_out1_valid}), .ready_out_bus({Buffer_15_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n5 (.clk(phi_n5_clk), .rst(phi_n5_rst), .data_in_bus({phi_n5_in2_data, phi_n5_in1_data}), .valid_in_bus({phi_n5_in2_valid, phi_n5_in1_valid}), .ready_in_bus({phi_n5_in2_ready, phi_n5_in1_ready}), .data_out_bus({phi_n5_out1_data}), .valid_out_bus({phi_n5_out1_valid}), .ready_out_bus({phi_n5_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_20 (.clk(fork_20_clk), .rst(fork_20_rst), .data_in_bus({fork_20_in1_data}), .valid_in_bus({fork_20_in1_valid}), .ready_in_bus({fork_20_in1_ready}), .data_out_bus({fork_20_out2_data, fork_20_out1_data}), .valid_out_bus({fork_20_out2_valid, fork_20_out1_valid}), .ready_out_bus({fork_20_out2_ready, fork_20_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_10 (.clk(source_10_clk), .rst(source_10_rst), .data_out_bus({source_10_out1_data}), .valid_out_bus({source_10_out1_valid}), .ready_out_bus({source_10_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_1 (.clk(branch_1_clk), .rst(branch_1_rst), .data_in_bus({{31'b0, branch_1_in2_data}, branch_1_in1_data}), .valid_in_bus({branch_1_in2_valid, branch_1_in1_valid}), .ready_in_bus({branch_1_in2_ready, branch_1_in1_ready}), .data_out_bus({branch_1_out2_data, branch_1_out1_data}), .valid_out_bus({branch_1_out2_valid, branch_1_out1_valid}), .ready_out_bus({branch_1_out2_ready, branch_1_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) OEHB_Buffer_25 (.clk(Buffer_25_clk), .rst(Buffer_25_rst), .data_in_bus({Buffer_25_in1_data}), .valid_in_bus({Buffer_25_in1_valid}), .ready_in_bus({Buffer_25_in1_ready}), .data_out_bus({Buffer_25_out1_data}), .valid_out_bus({Buffer_25_out1_valid}), .ready_out_bus({Buffer_25_out1_ready}));
mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_82 (.clk(phi_82_clk), .rst(phi_82_rst), .data_in_bus({{31'b0, phi_82_in1_data}, phi_82_in3_data, phi_82_in2_data}), .valid_in_bus({phi_82_in1_valid, phi_82_in3_valid, phi_82_in2_valid}), .ready_in_bus({phi_82_in1_ready, phi_82_in3_ready, phi_82_in2_ready}), .data_out_bus({phi_82_out1_data}), .valid_out_bus({phi_82_out1_valid}), .ready_out_bus({phi_82_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_1 (.clk(Buffer_1_clk), .rst(Buffer_1_rst), .data_in_bus({Buffer_1_in1_data}), .valid_in_bus({Buffer_1_in1_valid}), .ready_in_bus({Buffer_1_in1_ready}), .data_out_bus({Buffer_1_out1_data}), .valid_out_bus({Buffer_1_out1_valid}), .ready_out_bus({Buffer_1_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_36 (.clk(sink_36_clk), .rst(sink_36_rst), .data_in_bus({sink_36_in1_data}), .valid_in_bus({sink_36_in1_valid}), .ready_in_bus({sink_36_in1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_16 (.clk(cst_16_clk), .rst(cst_16_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_16_in1_valid}), .ready_in_bus({cst_16_in1_ready}), .data_out_bus({cst_16_out1_data}), .valid_out_bus({cst_16_out1_valid}), .ready_out_bus({cst_16_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_32 (.clk(fork_32_clk), .rst(fork_32_rst), .data_in_bus({fork_32_in1_data}), .valid_in_bus({fork_32_in1_valid}), .ready_in_bus({fork_32_in1_ready}), .data_out_bus({fork_32_out4_data, fork_32_out3_data, fork_32_out2_data, fork_32_out1_data}), .valid_out_bus({fork_32_out4_valid, fork_32_out3_valid, fork_32_out2_valid, fork_32_out1_valid}), .ready_out_bus({fork_32_out4_ready, fork_32_out3_ready, fork_32_out2_ready, fork_32_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_13 (.clk(branch_13_clk), .rst(branch_13_rst), .data_in_bus({{31'b0, branch_13_in2_data}, branch_13_in1_data}), .valid_in_bus({branch_13_in2_valid, branch_13_in1_valid}), .ready_in_bus({branch_13_in2_ready, branch_13_in1_ready}), .data_out_bus({branch_13_out2_data, branch_13_out1_data}), .valid_out_bus({branch_13_out2_valid, branch_13_out1_valid}), .ready_out_bus({branch_13_out2_ready, branch_13_out1_ready}));
MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(2), .LOAD_COUNT(3), .STORE_COUNT(2))MemCont_MC_x (.clk(MC_x_clk), .rst(MC_x_rst), .io_storeDataOut(x_dout0), .io_storeAddrOut(x_address0), .io_storeEnable(x_we0), .io_loadDataIn(x_din1), .io_loadAddrOut(x_address1), .io_loadEnable(x_ce1), .io_bbpValids({MC_x_in2_valid, MC_x_in1_valid}), .io_bb_stCountArray({MC_x_in2_data, MC_x_in1_data}), .io_bbReadyToPrevs({MC_x_in2_ready, MC_x_in1_ready}), .io_rdPortsPrev_ready({MC_x_in9_ready, MC_x_in6_ready, MC_x_in3_ready}), .io_rdPortsPrev_valid({MC_x_in9_valid, MC_x_in6_valid, MC_x_in3_valid}), .io_rdPortsPrev_bits({MC_x_in9_data, MC_x_in6_data, MC_x_in3_data}), .io_wrAddrPorts_ready({MC_x_in7_ready, MC_x_in4_ready}), .io_wrAddrPorts_valid({MC_x_in7_valid, MC_x_in4_valid}), .io_wrAddrPorts_bits({MC_x_in7_data, MC_x_in4_data}), .io_wrDataPorts_ready({MC_x_in8_ready, MC_x_in5_ready}), .io_wrDataPorts_valid({MC_x_in8_valid, MC_x_in5_valid}), .io_wrDataPorts_bits({MC_x_in8_data, MC_x_in5_data}), .io_rdPortsNext_ready({MC_x_out3_ready, MC_x_out2_ready, MC_x_out1_ready}), .io_rdPortsNext_valid({MC_x_out3_valid, MC_x_out2_valid, MC_x_out1_valid}), .io_rdPortsNext_bits({MC_x_out3_data, MC_x_out2_data, MC_x_out1_data}), .io_Empty_Valid({MC_x_out4_valid}), .io_Empty_Ready({MC_x_out4_ready}));
shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(11), .DATA_OUT_SIZE(11)) shl_op_shl_25 (.clk(shl_25_clk), .rst(shl_25_rst), .data_in_bus({shl_25_in2_data, shl_25_in1_data}), .valid_in_bus({shl_25_in2_valid, shl_25_in1_valid}), .ready_in_bus({shl_25_in2_ready, shl_25_in1_ready}), .data_out_bus({shl_25_out1_data}), .valid_out_bus({shl_25_out1_valid}), .ready_out_bus({shl_25_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_100 (.clk(add_100_clk), .rst(add_100_rst), .data_in_bus({add_100_in2_data, add_100_in1_data}), .valid_in_bus({add_100_in2_valid, add_100_in1_valid}), .ready_in_bus({add_100_in2_ready, add_100_in1_ready}), .data_out_bus({add_100_out1_data}), .valid_out_bus({add_100_out1_valid}), .ready_out_bus({add_100_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_22 (.clk(sink_22_clk), .rst(sink_22_rst), .data_in_bus({sink_22_in1_data}), .valid_in_bus({sink_22_in1_valid}), .ready_in_bus({sink_22_in1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_14 (.clk(source_14_clk), .rst(source_14_rst), .data_out_bus({source_14_out1_data}), .valid_out_bus({source_14_out1_valid}), .ready_out_bus({source_14_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) OEHB_Buffer_2 (.clk(Buffer_2_clk), .rst(Buffer_2_rst), .data_in_bus({Buffer_2_in1_data}), .valid_in_bus({Buffer_2_in1_valid}), .ready_in_bus({Buffer_2_in1_ready}), .data_out_bus({Buffer_2_out1_data}), .valid_out_bus({Buffer_2_out1_valid}), .ready_out_bus({Buffer_2_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_15 (.clk(sink_15_clk), .rst(sink_15_rst), .data_in_bus({sink_15_in1_data}), .valid_in_bus({sink_15_in1_valid}), .ready_in_bus({sink_15_in1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n26 (.clk(phi_n26_clk), .rst(phi_n26_rst), .data_in_bus({phi_n26_in2_data, phi_n26_in1_data}), .valid_in_bus({phi_n26_in2_valid, phi_n26_in1_valid}), .ready_in_bus({phi_n26_in2_ready, phi_n26_in1_ready}), .data_out_bus({phi_n26_out1_data}), .valid_out_bus({phi_n26_out1_valid}), .ready_out_bus({phi_n26_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_12 (.clk(source_12_clk), .rst(source_12_rst), .data_out_bus({source_12_out1_data}), .valid_out_bus({source_12_out1_valid}), .ready_out_bus({source_12_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(12), .DATA_SIZE(32)) mc_load_op_load_88 (.clk(load_88_clk), .rst(load_88_rst), .data_in_bus({load_88_in1_data}), .address_in_bus({load_88_in2_data}), .valid_in_bus({load_88_in2_valid, load_88_in1_valid}), .ready_in_bus({load_88_in2_ready, load_88_in1_ready}), .data_out_bus({load_88_out1_data}), .address_out_bus({load_88_out2_data}), .valid_out_bus({load_88_out2_valid, load_88_out1_valid}), .ready_out_bus({load_88_out2_ready, load_88_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_17 (.clk(source_17_clk), .rst(source_17_rst), .data_out_bus({source_17_out1_data}), .valid_out_bus({source_17_out1_valid}), .ready_out_bus({source_17_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n19 (.clk(phi_n19_clk), .rst(phi_n19_rst), .data_in_bus({phi_n19_in1_data}), .valid_in_bus({phi_n19_in1_valid}), .ready_in_bus({phi_n19_in1_ready}), .data_out_bus({phi_n19_out1_data}), .valid_out_bus({phi_n19_out1_valid}), .ready_out_bus({phi_n19_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_32 (.clk(sink_32_clk), .rst(sink_32_rst), .data_in_bus({sink_32_in1_data}), .valid_in_bus({sink_32_in1_valid}), .ready_in_bus({sink_32_in1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_6 (.clk(fork_6_clk), .rst(fork_6_rst), .data_in_bus({fork_6_in1_data}), .valid_in_bus({fork_6_in1_valid}), .ready_in_bus({fork_6_in1_ready}), .data_out_bus({fork_6_out2_data, fork_6_out1_data}), .valid_out_bus({fork_6_out2_valid, fork_6_out1_valid}), .ready_out_bus({fork_6_out2_ready, fork_6_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_15 (.clk(source_15_clk), .rst(source_15_rst), .data_out_bus({source_15_out1_data}), .valid_out_bus({source_15_out1_valid}), .ready_out_bus({source_15_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_16 (.clk(add_16_clk), .rst(add_16_rst), .data_in_bus({add_16_in2_data, add_16_in1_data}), .valid_in_bus({add_16_in2_valid, add_16_in1_valid}), .ready_in_bus({add_16_in2_ready, add_16_in1_ready}), .data_out_bus({add_16_out1_data}), .valid_out_bus({add_16_out1_valid}), .ready_out_bus({add_16_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_8 (.clk(source_8_clk), .rst(source_8_rst), .data_out_bus({source_8_out1_data}), .valid_out_bus({source_8_out1_valid}), .ready_out_bus({source_8_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_11 (.clk(load_11_clk), .rst(load_11_rst), .data_in_bus({load_11_in1_data}), .address_in_bus({load_11_in2_data}), .valid_in_bus({load_11_in2_valid, load_11_in1_valid}), .ready_in_bus({load_11_in2_ready, load_11_in1_ready}), .data_out_bus({load_11_out1_data}), .address_out_bus({load_11_out2_data}), .valid_out_bus({load_11_out2_valid, load_11_out1_valid}), .ready_out_bus({load_11_out2_ready, load_11_out1_ready}));
start_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) start_node_alpha (.clk(alpha_clk), .rst(alpha_rst), .data_in_bus({alpha_in1_data}), .valid_in_bus({alpha_in1_valid}), .ready_in_bus({alpha_in1_ready}), .data_out_bus({alpha_out1_data}), .valid_out_bus({alpha_out1_valid}), .ready_out_bus({alpha_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_73 (.clk(add_73_clk), .rst(add_73_rst), .data_in_bus({add_73_in2_data, add_73_in1_data}), .valid_in_bus({add_73_in2_valid, add_73_in1_valid}), .ready_in_bus({add_73_in2_ready, add_73_in1_ready}), .data_out_bus({add_73_out1_data}), .valid_out_bus({add_73_out1_valid}), .ready_out_bus({add_73_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_4 (.clk(source_4_clk), .rst(source_4_rst), .data_out_bus({source_4_out1_data}), .valid_out_bus({source_4_out1_valid}), .ready_out_bus({source_4_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_54 (.clk(add_54_clk), .rst(add_54_rst), .data_in_bus({add_54_in2_data, add_54_in1_data}), .valid_in_bus({add_54_in2_valid, add_54_in1_valid}), .ready_in_bus({add_54_in2_ready, add_54_in1_ready}), .data_out_bus({add_54_out1_data}), .valid_out_bus({add_54_out1_valid}), .ready_out_bus({add_54_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_9 (.clk(source_9_clk), .rst(source_9_rst), .data_out_bus({source_9_out1_data}), .valid_out_bus({source_9_out1_valid}), .ready_out_bus({source_9_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_37 (.clk(branch_37_clk), .rst(branch_37_rst), .data_in_bus({{branch_37_in2_data}, branch_37_in1_data}), .valid_in_bus({branch_37_in2_valid, branch_37_in1_valid}), .ready_in_bus({branch_37_in2_ready, branch_37_in1_ready}), .data_out_bus({branch_37_out2_data, branch_37_out1_data}), .valid_out_bus({branch_37_out2_valid, branch_37_out1_valid}), .ready_out_bus({branch_37_out2_ready, branch_37_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_37 (.clk(phiC_37_clk), .rst(phiC_37_rst), .data_in_bus({phiC_37_in1_data}), .valid_in_bus({phiC_37_in1_valid}), .ready_in_bus({phiC_37_in1_ready}), .data_out_bus({phiC_37_out1_data}), .valid_out_bus({phiC_37_out1_valid}), .ready_out_bus({phiC_37_out1_ready}));
MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_v1 (.clk(MC_v1_clk), .rst(MC_v1_rst), .io_storeDataOut(v1_dout0), .io_storeAddrOut(v1_address0), .io_storeEnable(v1_we0), .io_loadDataIn(v1_din1), .io_loadAddrOut(v1_address1), .io_loadEnable(v1_ce1), .io_bbpValids({MC_v1_in2_valid}), .io_bb_stCountArray({MC_v1_in2_data}), .io_bbReadyToPrevs({MC_v1_in2_ready}), .io_rdPortsPrev_ready({MC_v1_in1_ready}), .io_rdPortsPrev_valid({MC_v1_in1_valid}), .io_rdPortsPrev_bits({MC_v1_in1_data}), .io_wrAddrPorts_ready({MC_v1_in3_ready}), .io_wrAddrPorts_valid({MC_v1_in3_valid}), .io_wrAddrPorts_bits({MC_v1_in3_data}), .io_wrDataPorts_ready({MC_v1_in4_ready}), .io_wrDataPorts_valid({MC_v1_in4_valid}), .io_wrDataPorts_bits({MC_v1_in4_data}), .io_rdPortsNext_ready({MC_v1_out1_ready}), .io_rdPortsNext_valid({MC_v1_out1_valid}), .io_rdPortsNext_bits({MC_v1_out1_data}), .io_Empty_Valid({MC_v1_out2_valid}), .io_Empty_Ready({MC_v1_out2_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_2 (.clk(cst_2_clk), .rst(cst_2_rst), .data_in_bus({3'd5}), .valid_in_bus({cst_2_in1_valid}), .ready_in_bus({cst_2_in1_ready}), .data_out_bus({cst_2_out1_data}), .valid_out_bus({cst_2_out1_valid}), .ready_out_bus({cst_2_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n18 (.clk(phi_n18_clk), .rst(phi_n18_rst), .data_in_bus({phi_n18_in2_data, phi_n18_in1_data}), .valid_in_bus({phi_n18_in2_valid, phi_n18_in1_valid}), .ready_in_bus({phi_n18_in2_ready, phi_n18_in1_ready}), .data_out_bus({phi_n18_out1_data}), .valid_out_bus({phi_n18_out1_valid}), .ready_out_bus({phi_n18_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_57 (.clk(branchC_57_clk), .rst(branchC_57_rst), .data_in_bus({{branchC_57_in2_data}, branchC_57_in1_data}), .valid_in_bus({branchC_57_in2_valid, branchC_57_in1_valid}), .ready_in_bus({branchC_57_in2_ready, branchC_57_in1_ready}), .data_out_bus({branchC_57_out2_data, branchC_57_out1_data}), .valid_out_bus({branchC_57_out2_valid, branchC_57_out1_valid}), .ready_out_bus({branchC_57_out2_ready, branchC_57_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_94 (.clk(add_94_clk), .rst(add_94_rst), .data_in_bus({add_94_in2_data, add_94_in1_data}), .valid_in_bus({add_94_in2_valid, add_94_in1_valid}), .ready_in_bus({add_94_in2_ready, add_94_in1_ready}), .data_out_bus({add_94_out1_data}), .valid_out_bus({add_94_out1_valid}), .ready_out_bus({add_94_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n16 (.clk(phi_n16_clk), .rst(phi_n16_rst), .data_in_bus({phi_n16_in2_data, phi_n16_in1_data}), .valid_in_bus({phi_n16_in2_valid, phi_n16_in1_valid}), .ready_in_bus({phi_n16_in2_ready, phi_n16_in1_ready}), .data_out_bus({phi_n16_out1_data}), .valid_out_bus({phi_n16_out1_valid}), .ready_out_bus({phi_n16_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_14 (.clk(load_14_clk), .rst(load_14_rst), .data_in_bus({load_14_in1_data}), .address_in_bus({load_14_in2_data}), .valid_in_bus({load_14_in2_valid, load_14_in1_valid}), .ready_in_bus({load_14_in2_ready, load_14_in1_ready}), .data_out_bus({load_14_out1_data}), .address_out_bus({load_14_out2_data}), .valid_out_bus({load_14_out2_valid, load_14_out1_valid}), .ready_out_bus({load_14_out2_ready, load_14_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_5 (.clk(branch_5_clk), .rst(branch_5_rst), .data_in_bus({{31'b0, branch_5_in2_data}, branch_5_in1_data}), .valid_in_bus({branch_5_in2_valid, branch_5_in1_valid}), .ready_in_bus({branch_5_in2_ready, branch_5_in1_ready}), .data_out_bus({branch_5_out2_data, branch_5_out1_data}), .valid_out_bus({branch_5_out2_valid, branch_5_out1_valid}), .ready_out_bus({branch_5_out2_ready, branch_5_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_11 (.clk(Buffer_11_clk), .rst(Buffer_11_rst), .data_in_bus({Buffer_11_in1_data}), .valid_in_bus({Buffer_11_in1_valid}), .ready_in_bus({Buffer_11_in1_ready}), .data_out_bus({Buffer_11_out1_data}), .valid_out_bus({Buffer_11_out1_valid}), .ready_out_bus({Buffer_11_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_19 (.clk(Buffer_19_clk), .rst(Buffer_19_rst), .data_in_bus({Buffer_19_in1_data}), .valid_in_bus({Buffer_19_in1_valid}), .ready_in_bus({Buffer_19_in1_ready}), .data_out_bus({Buffer_19_out1_data}), .valid_out_bus({Buffer_19_out1_valid}), .ready_out_bus({Buffer_19_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_8 (.clk(Buffer_8_clk), .rst(Buffer_8_rst), .data_in_bus({Buffer_8_in1_data}), .valid_in_bus({Buffer_8_in1_valid}), .ready_in_bus({Buffer_8_in1_ready}), .data_out_bus({Buffer_8_out1_data}), .valid_out_bus({Buffer_8_out1_valid}), .ready_out_bus({Buffer_8_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_23 (.clk(Buffer_23_clk), .rst(Buffer_23_rst), .data_in_bus({Buffer_23_in1_data}), .valid_in_bus({Buffer_23_in1_valid}), .ready_in_bus({Buffer_23_in1_ready}), .data_out_bus({Buffer_23_out1_data}), .valid_out_bus({Buffer_23_out1_valid}), .ready_out_bus({Buffer_23_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_33 (.clk(fork_33_clk), .rst(fork_33_rst), .data_in_bus({fork_33_in1_data}), .valid_in_bus({fork_33_in1_valid}), .ready_in_bus({fork_33_in1_ready}), .data_out_bus({fork_33_out4_data, fork_33_out3_data, fork_33_out2_data, fork_33_out1_data}), .valid_out_bus({fork_33_out4_valid, fork_33_out3_valid, fork_33_out2_valid, fork_33_out1_valid}), .ready_out_bus({fork_33_out4_ready, fork_33_out3_ready, fork_33_out2_ready, fork_33_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_29 (.clk(add_29_clk), .rst(add_29_rst), .data_in_bus({add_29_in2_data, add_29_in1_data}), .valid_in_bus({add_29_in2_valid, add_29_in1_valid}), .ready_in_bus({add_29_in2_ready, add_29_in1_ready}), .data_out_bus({add_29_out1_data}), .valid_out_bus({add_29_out1_valid}), .ready_out_bus({add_29_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_51 (.clk(forkC_51_clk), .rst(forkC_51_rst), .data_in_bus({forkC_51_in1_data}), .valid_in_bus({forkC_51_in1_valid}), .ready_in_bus({forkC_51_in1_ready}), .data_out_bus({forkC_51_out2_data, forkC_51_out1_data}), .valid_out_bus({forkC_51_out2_valid, forkC_51_out1_valid}), .ready_out_bus({forkC_51_out2_ready, forkC_51_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_31 (.clk(sink_31_clk), .rst(sink_31_rst), .data_in_bus({sink_31_in1_data}), .valid_in_bus({sink_31_in1_valid}), .ready_in_bus({sink_31_in1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) OEHB_Buffer_0 (.clk(Buffer_0_clk), .rst(Buffer_0_rst), .data_in_bus({Buffer_0_in1_data}), .valid_in_bus({Buffer_0_in1_valid}), .ready_in_bus({Buffer_0_in1_ready}), .data_out_bus({Buffer_0_out1_data}), .valid_out_bus({Buffer_0_out1_valid}), .ready_out_bus({Buffer_0_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_27 (.clk(cst_27_clk), .rst(cst_27_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_27_in1_valid}), .ready_in_bus({cst_27_in1_ready}), .data_out_bus({cst_27_out1_data}), .valid_out_bus({cst_27_out1_valid}), .ready_out_bus({cst_27_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_19 (.clk(load_19_clk), .rst(load_19_rst), .data_in_bus({load_19_in1_data}), .address_in_bus({load_19_in2_data}), .valid_in_bus({load_19_in2_valid, load_19_in1_valid}), .ready_in_bus({load_19_in2_ready, load_19_in1_ready}), .data_out_bus({load_19_out1_data}), .address_out_bus({load_19_out2_data}), .valid_out_bus({load_19_out2_valid, load_19_out1_valid}), .ready_out_bus({load_19_out2_ready, load_19_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n20 (.clk(phi_n20_clk), .rst(phi_n20_rst), .data_in_bus({phi_n20_in2_data, phi_n20_in1_data}), .valid_in_bus({phi_n20_in2_valid, phi_n20_in1_valid}), .ready_in_bus({phi_n20_in2_ready, phi_n20_in1_ready}), .data_out_bus({phi_n20_out1_data}), .valid_out_bus({phi_n20_out1_valid}), .ready_out_bus({phi_n20_out1_ready}));
icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_74 (.clk(icmp_74_clk), .rst(icmp_74_rst), .data_in_bus({icmp_74_in2_data, icmp_74_in1_data}), .valid_in_bus({icmp_74_in2_valid, icmp_74_in1_valid}), .ready_in_bus({icmp_74_in2_ready, icmp_74_in1_ready}), .data_out_bus({icmp_74_out1_data}), .valid_out_bus({icmp_74_out1_valid}), .ready_out_bus({icmp_74_out1_ready}));
shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(11), .DATA_OUT_SIZE(11)) shl_op_shl_4 (.clk(shl_4_clk), .rst(shl_4_rst), .data_in_bus({shl_4_in2_data, shl_4_in1_data}), .valid_in_bus({shl_4_in2_valid, shl_4_in1_valid}), .ready_in_bus({shl_4_in2_ready, shl_4_in1_ready}), .data_out_bus({shl_4_out1_data}), .valid_out_bus({shl_4_out1_valid}), .ready_out_bus({shl_4_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_4 (.clk(branch_4_clk), .rst(branch_4_rst), .data_in_bus({{5'b0, branch_4_in2_data}, branch_4_in1_data}), .valid_in_bus({branch_4_in2_valid, branch_4_in1_valid}), .ready_in_bus({branch_4_in2_ready, branch_4_in1_ready}), .data_out_bus({branch_4_out2_data, branch_4_out1_data}), .valid_out_bus({branch_4_out2_valid, branch_4_out1_valid}), .ready_out_bus({branch_4_out2_ready, branch_4_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n2 (.clk(phi_n2_clk), .rst(phi_n2_rst), .data_in_bus({phi_n2_in1_data}), .valid_in_bus({phi_n2_in1_valid}), .ready_in_bus({phi_n2_in1_ready}), .data_out_bus({phi_n2_out1_data}), .valid_out_bus({phi_n2_out1_valid}), .ready_out_bus({phi_n2_out1_ready}));
mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_77 (.clk(phi_77_clk), .rst(phi_77_rst), .data_in_bus({{5'b0, phi_77_in1_data}, phi_77_in3_data, phi_77_in2_data}), .valid_in_bus({phi_77_in1_valid, phi_77_in3_valid, phi_77_in2_valid}), .ready_in_bus({phi_77_in1_ready, phi_77_in3_ready, phi_77_in2_ready}), .data_out_bus({phi_77_out1_data}), .valid_out_bus({phi_77_out1_valid}), .ready_out_bus({phi_77_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_47 (.clk(branchC_47_clk), .rst(branchC_47_rst), .data_in_bus({{branchC_47_in2_data}, branchC_47_in1_data}), .valid_in_bus({branchC_47_in2_valid, branchC_47_in1_valid}), .ready_in_bus({branchC_47_in2_ready, branchC_47_in1_ready}), .data_out_bus({branchC_47_out2_data, branchC_47_out1_data}), .valid_out_bus({branchC_47_out2_valid, branchC_47_out1_valid}), .ready_out_bus({branchC_47_out2_ready, branchC_47_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_44 (.clk(branch_44_clk), .rst(branch_44_rst), .data_in_bus({{31'b0, branch_44_in2_data}, branch_44_in1_data}), .valid_in_bus({branch_44_in2_valid, branch_44_in1_valid}), .ready_in_bus({branch_44_in2_ready, branch_44_in1_ready}), .data_out_bus({branch_44_out2_data, branch_44_out1_data}), .valid_out_bus({branch_44_out2_valid, branch_44_out1_valid}), .ready_out_bus({branch_44_out2_ready, branch_44_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_29 (.clk(fork_29_clk), .rst(fork_29_rst), .data_in_bus({fork_29_in1_data}), .valid_in_bus({fork_29_in1_valid}), .ready_in_bus({fork_29_in1_ready}), .data_out_bus({fork_29_out4_data, fork_29_out3_data, fork_29_out2_data, fork_29_out1_data}), .valid_out_bus({fork_29_out4_valid, fork_29_out3_valid, fork_29_out2_valid, fork_29_out1_valid}), .ready_out_bus({fork_29_out4_ready, fork_29_out3_ready, fork_29_out2_ready, fork_29_out1_ready}));
MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_u1 (.clk(MC_u1_clk), .rst(MC_u1_rst), .io_storeDataOut(u1_dout0), .io_storeAddrOut(u1_address0), .io_storeEnable(u1_we0), .io_loadDataIn(u1_din1), .io_loadAddrOut(u1_address1), .io_loadEnable(u1_ce1), .io_bbpValids({MC_u1_in2_valid}), .io_bb_stCountArray({MC_u1_in2_data}), .io_bbReadyToPrevs({MC_u1_in2_ready}), .io_rdPortsPrev_ready({MC_u1_in1_ready}), .io_rdPortsPrev_valid({MC_u1_in1_valid}), .io_rdPortsPrev_bits({MC_u1_in1_data}), .io_wrAddrPorts_ready({MC_u1_in3_ready}), .io_wrAddrPorts_valid({MC_u1_in3_valid}), .io_wrAddrPorts_bits({MC_u1_in3_data}), .io_wrDataPorts_ready({MC_u1_in4_ready}), .io_wrDataPorts_valid({MC_u1_in4_valid}), .io_wrDataPorts_bits({MC_u1_in4_data}), .io_rdPortsNext_ready({MC_u1_out1_ready}), .io_rdPortsNext_valid({MC_u1_out1_valid}), .io_rdPortsNext_bits({MC_u1_out1_data}), .io_Empty_Valid({MC_u1_out2_valid}), .io_Empty_Ready({MC_u1_out2_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_49 (.clk(forkC_49_clk), .rst(forkC_49_rst), .data_in_bus({forkC_49_in1_data}), .valid_in_bus({forkC_49_in1_valid}), .ready_in_bus({forkC_49_in1_ready}), .data_out_bus({forkC_49_out3_data, forkC_49_out2_data, forkC_49_out1_data}), .valid_out_bus({forkC_49_out3_valid, forkC_49_out2_valid, forkC_49_out1_valid}), .ready_out_bus({forkC_49_out3_ready, forkC_49_out2_ready, forkC_49_out1_ready}));
MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(12), .BB_COUNT(1), .LOAD_COUNT(3), .STORE_COUNT(1))MemCont_MC_A (.clk(MC_A_clk), .rst(MC_A_rst), .io_storeDataOut(A_dout0), .io_storeAddrOut(A_address0), .io_storeEnable(A_we0), .io_loadDataIn(A_din1), .io_loadAddrOut(A_address1), .io_loadEnable(A_ce1), .io_bbpValids({MC_A_in1_valid}), .io_bb_stCountArray({MC_A_in1_data}), .io_bbReadyToPrevs({MC_A_in1_ready}), .io_rdPortsPrev_ready({MC_A_in6_ready, MC_A_in5_ready, MC_A_in2_ready}), .io_rdPortsPrev_valid({MC_A_in6_valid, MC_A_in5_valid, MC_A_in2_valid}), .io_rdPortsPrev_bits({MC_A_in6_data, MC_A_in5_data, MC_A_in2_data}), .io_wrAddrPorts_ready({MC_A_in3_ready}), .io_wrAddrPorts_valid({MC_A_in3_valid}), .io_wrAddrPorts_bits({MC_A_in3_data}), .io_wrDataPorts_ready({MC_A_in4_ready}), .io_wrDataPorts_valid({MC_A_in4_valid}), .io_wrDataPorts_bits({MC_A_in4_data}), .io_rdPortsNext_ready({MC_A_out3_ready, MC_A_out2_ready, MC_A_out1_ready}), .io_rdPortsNext_valid({MC_A_out3_valid, MC_A_out2_valid, MC_A_out1_valid}), .io_rdPortsNext_bits({MC_A_out3_data, MC_A_out2_data, MC_A_out1_data}), .io_Empty_Valid({MC_A_out4_valid}), .io_Empty_Ready({MC_A_out4_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_23 (.clk(sink_23_clk), .rst(sink_23_rst), .data_in_bus({sink_23_in1_data}), .valid_in_bus({sink_23_in1_valid}), .ready_in_bus({sink_23_in1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_3 (.clk(fork_3_clk), .rst(fork_3_rst), .data_in_bus({fork_3_in1_data}), .valid_in_bus({fork_3_in1_valid}), .ready_in_bus({fork_3_in1_ready}), .data_out_bus({fork_3_out2_data, fork_3_out1_data}), .valid_out_bus({fork_3_out2_valid, fork_3_out1_valid}), .ready_out_bus({fork_3_out2_ready, fork_3_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_2 (.clk(sink_2_clk), .rst(sink_2_rst), .data_in_bus({sink_2_in1_data}), .valid_in_bus({sink_2_in1_valid}), .ready_in_bus({sink_2_in1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_34 (.clk(phiC_34_clk), .rst(phiC_34_rst), .data_in_bus({phiC_34_in1_data}), .valid_in_bus({phiC_34_in1_valid}), .ready_in_bus({phiC_34_in1_ready}), .data_out_bus({phiC_34_out1_data}), .valid_out_bus({phiC_34_out1_valid}), .ready_out_bus({phiC_34_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_12 (.clk(cst_12_clk), .rst(cst_12_rst), .data_in_bus({6'd32}), .valid_in_bus({cst_12_in1_valid}), .ready_in_bus({cst_12_in1_ready}), .data_out_bus({cst_12_out1_data}), .valid_out_bus({cst_12_out1_valid}), .ready_out_bus({cst_12_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_30 (.clk(sink_30_clk), .rst(sink_30_rst), .data_in_bus({sink_30_in1_data}), .valid_in_bus({sink_30_in1_valid}), .ready_in_bus({sink_30_in1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n1 (.clk(phi_n1_clk), .rst(phi_n1_rst), .data_in_bus({phi_n1_in2_data, phi_n1_in1_data}), .valid_in_bus({phi_n1_in2_valid, phi_n1_in1_valid}), .ready_in_bus({phi_n1_in2_ready, phi_n1_in1_ready}), .data_out_bus({phi_n1_out1_data}), .valid_out_bus({phi_n1_out1_valid}), .ready_out_bus({phi_n1_out1_ready}));
ret_op #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) ret_op_ret_0 (.clk(ret_0_clk), .rst(ret_0_rst), .data_in_bus({ret_0_in1_data}), .valid_in_bus({ret_0_in1_valid}), .ready_in_bus({ret_0_in1_ready}), .data_out_bus({ret_0_out1_data}), .valid_out_bus({ret_0_out1_valid}), .ready_out_bus({ret_0_out1_ready}));
mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_83 (.clk(phi_83_clk), .rst(phi_83_rst), .data_in_bus({{5'b0, phi_83_in1_data}, phi_83_in3_data, phi_83_in2_data}), .valid_in_bus({phi_83_in1_valid, phi_83_in3_valid, phi_83_in2_valid}), .ready_in_bus({phi_83_in1_ready, phi_83_in3_ready, phi_83_in2_ready}), .data_out_bus({phi_83_out1_data}), .valid_out_bus({phi_83_out1_valid}), .ready_out_bus({phi_83_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_66 (.clk(load_66_clk), .rst(load_66_rst), .data_in_bus({load_66_in1_data}), .address_in_bus({load_66_in2_data}), .valid_in_bus({load_66_in2_valid, load_66_in1_valid}), .ready_in_bus({load_66_in2_ready, load_66_in1_ready}), .data_out_bus({load_66_out1_data}), .address_out_bus({load_66_out2_data}), .valid_out_bus({load_66_out2_valid, load_66_out1_valid}), .ready_out_bus({load_66_out2_ready, load_66_out1_ready}));
MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_v2 (.clk(MC_v2_clk), .rst(MC_v2_rst), .io_storeDataOut(v2_dout0), .io_storeAddrOut(v2_address0), .io_storeEnable(v2_we0), .io_loadDataIn(v2_din1), .io_loadAddrOut(v2_address1), .io_loadEnable(v2_ce1), .io_bbpValids({MC_v2_in2_valid}), .io_bb_stCountArray({MC_v2_in2_data}), .io_bbReadyToPrevs({MC_v2_in2_ready}), .io_rdPortsPrev_ready({MC_v2_in1_ready}), .io_rdPortsPrev_valid({MC_v2_in1_valid}), .io_rdPortsPrev_bits({MC_v2_in1_data}), .io_wrAddrPorts_ready({MC_v2_in3_ready}), .io_wrAddrPorts_valid({MC_v2_in3_valid}), .io_wrAddrPorts_bits({MC_v2_in3_data}), .io_wrDataPorts_ready({MC_v2_in4_ready}), .io_wrDataPorts_valid({MC_v2_in4_valid}), .io_wrDataPorts_bits({MC_v2_in4_data}), .io_rdPortsNext_ready({MC_v2_out1_ready}), .io_rdPortsNext_valid({MC_v2_out1_valid}), .io_rdPortsNext_bits({MC_v2_out1_data}), .io_Empty_Valid({MC_v2_out2_valid}), .io_Empty_Ready({MC_v2_out2_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_20 (.clk(sink_20_clk), .rst(sink_20_rst), .data_in_bus({sink_20_in1_data}), .valid_in_bus({sink_20_in1_valid}), .ready_in_bus({sink_20_in1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) OEHB_Buffer_26 (.clk(Buffer_26_clk), .rst(Buffer_26_rst), .data_in_bus({Buffer_26_in1_data}), .valid_in_bus({Buffer_26_in1_valid}), .ready_in_bus({Buffer_26_in1_ready}), .data_out_bus({Buffer_26_out1_data}), .valid_out_bus({Buffer_26_out1_valid}), .ready_out_bus({Buffer_26_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_26 (.clk(branch_26_clk), .rst(branch_26_rst), .data_in_bus({{31'b0, branch_26_in2_data}, branch_26_in1_data}), .valid_in_bus({branch_26_in2_valid, branch_26_in1_valid}), .ready_in_bus({branch_26_in2_ready, branch_26_in1_ready}), .data_out_bus({branch_26_out2_data, branch_26_out1_data}), .valid_out_bus({branch_26_out2_valid, branch_26_out1_valid}), .ready_out_bus({branch_26_out2_ready, branch_26_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_13 (.clk(cst_13_clk), .rst(cst_13_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_13_in1_valid}), .ready_in_bus({cst_13_in1_ready}), .data_out_bus({cst_13_out1_data}), .valid_out_bus({cst_13_out1_valid}), .ready_out_bus({cst_13_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_39 (.clk(branch_39_clk), .rst(branch_39_rst), .data_in_bus({{5'b0, branch_39_in2_data}, branch_39_in1_data}), .valid_in_bus({branch_39_in2_valid, branch_39_in1_valid}), .ready_in_bus({branch_39_in2_ready, branch_39_in1_ready}), .data_out_bus({branch_39_out2_data, branch_39_out1_data}), .valid_out_bus({branch_39_out2_valid, branch_39_out1_valid}), .ready_out_bus({branch_39_out2_ready, branch_39_out1_ready}));
mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(16), .DATA_OUT_SIZE(32)) mul_op_mul_89 (.clk(mul_89_clk), .rst(mul_89_rst), .data_in_bus({mul_89_in2_data, mul_89_in1_data}), .valid_in_bus({mul_89_in2_valid, mul_89_in1_valid}), .ready_in_bus({mul_89_in2_ready, mul_89_in1_ready}), .data_out_bus({mul_89_out1_data}), .valid_out_bus({mul_89_out1_valid}), .ready_out_bus({mul_89_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block6 (.clk(brCst_block6_clk), .rst(brCst_block6_rst), .data_in_bus({1'd1}), .valid_in_bus({brCst_block6_in1_valid}), .ready_in_bus({brCst_block6_in1_ready}), .data_out_bus({brCst_block6_out1_data}), .valid_out_bus({brCst_block6_out1_valid}), .ready_out_bus({brCst_block6_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_8 (.clk(branch_8_clk), .rst(branch_8_rst), .data_in_bus({{5'b0, branch_8_in2_data}, branch_8_in1_data}), .valid_in_bus({branch_8_in2_valid, branch_8_in1_valid}), .ready_in_bus({branch_8_in2_ready, branch_8_in1_ready}), .data_out_bus({branch_8_out2_data, branch_8_out1_data}), .valid_out_bus({branch_8_out2_valid, branch_8_out1_valid}), .ready_out_bus({branch_8_out2_ready, branch_8_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_51 (.clk(load_51_clk), .rst(load_51_rst), .data_in_bus({load_51_in1_data}), .address_in_bus({load_51_in2_data}), .valid_in_bus({load_51_in2_valid, load_51_in1_valid}), .ready_in_bus({load_51_in2_ready, load_51_in1_ready}), .data_out_bus({load_51_out1_data}), .address_out_bus({load_51_out2_data}), .valid_out_bus({load_51_out2_valid, load_51_out1_valid}), .ready_out_bus({load_51_out2_ready, load_51_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_0 (.clk(fork_0_clk), .rst(fork_0_rst), .data_in_bus({fork_0_in1_data}), .valid_in_bus({fork_0_in1_valid}), .ready_in_bus({fork_0_in1_ready}), .data_out_bus({fork_0_out5_data, fork_0_out4_data, fork_0_out3_data, fork_0_out2_data, fork_0_out1_data}), .valid_out_bus({fork_0_out5_valid, fork_0_out4_valid, fork_0_out3_valid, fork_0_out2_valid, fork_0_out1_valid}), .ready_out_bus({fork_0_out5_ready, fork_0_out4_ready, fork_0_out3_ready, fork_0_out2_ready, fork_0_out1_ready}));
mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_store_op_store_2 (.clk(store_2_clk), .rst(store_2_rst), .data_in_bus({store_2_in1_data}), .address_in_bus({store_2_in2_data}), .valid_in_bus({store_2_in2_valid, store_2_in1_valid}), .ready_in_bus({store_2_in2_ready, store_2_in1_ready}), .data_out_bus({store_2_out1_data}), .address_out_bus({store_2_out2_data}), .valid_out_bus({store_2_out2_valid, store_2_out1_valid}), .ready_out_bus({store_2_out2_ready, store_2_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_0 (.clk(cst_0_clk), .rst(cst_0_rst), .data_in_bus({1'd0}), .valid_in_bus({cst_0_in1_valid}), .ready_in_bus({cst_0_in1_ready}), .data_out_bus({cst_0_out1_data}), .valid_out_bus({cst_0_out1_valid}), .ready_out_bus({cst_0_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_14 (.clk(branch_14_clk), .rst(branch_14_rst), .data_in_bus({{branch_14_in2_data}, branch_14_in1_data}), .valid_in_bus({branch_14_in2_valid, branch_14_in1_valid}), .ready_in_bus({branch_14_in2_ready, branch_14_in1_ready}), .data_out_bus({branch_14_out2_data, branch_14_out1_data}), .valid_out_bus({branch_14_out2_valid, branch_14_out1_valid}), .ready_out_bus({branch_14_out2_ready, branch_14_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_58 (.clk(branchC_58_clk), .rst(branchC_58_rst), .data_in_bus({{branchC_58_in2_data}, branchC_58_in1_data}), .valid_in_bus({branchC_58_in2_valid, branchC_58_in1_valid}), .ready_in_bus({branchC_58_in2_ready, branchC_58_in1_ready}), .data_out_bus({branchC_58_out2_data, branchC_58_out1_data}), .valid_out_bus({branchC_58_out2_valid, branchC_58_out1_valid}), .ready_out_bus({branchC_58_out2_ready, branchC_58_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_3 (.clk(cst_3_clk), .rst(cst_3_rst), .data_in_bus({3'd5}), .valid_in_bus({cst_3_in1_valid}), .ready_in_bus({cst_3_in1_ready}), .data_out_bus({cst_3_out1_data}), .valid_out_bus({cst_3_out1_valid}), .ready_out_bus({cst_3_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_1 (.clk(cst_1_clk), .rst(cst_1_rst), .data_in_bus({1'd0}), .valid_in_bus({cst_1_in1_valid}), .ready_in_bus({cst_1_in1_ready}), .data_out_bus({cst_1_out1_data}), .valid_out_bus({cst_1_out1_valid}), .ready_out_bus({cst_1_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_0 (.clk(branch_0_clk), .rst(branch_0_rst), .data_in_bus({{branch_0_in2_data}, branch_0_in1_data}), .valid_in_bus({branch_0_in2_valid, branch_0_in1_valid}), .ready_in_bus({branch_0_in2_ready, branch_0_in1_ready}), .data_out_bus({branch_0_out2_data, branch_0_out1_data}), .valid_out_bus({branch_0_out2_valid, branch_0_out1_valid}), .ready_out_bus({branch_0_out2_ready, branch_0_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_28 (.clk(cst_28_clk), .rst(cst_28_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_28_in1_valid}), .ready_in_bus({cst_28_in1_ready}), .data_out_bus({cst_28_out1_data}), .valid_out_bus({cst_28_out1_valid}), .ready_out_bus({cst_28_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(6), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_34 (.clk(fork_34_clk), .rst(fork_34_rst), .data_in_bus({fork_34_in1_data}), .valid_in_bus({fork_34_in1_valid}), .ready_in_bus({fork_34_in1_ready}), .data_out_bus({fork_34_out6_data, fork_34_out5_data, fork_34_out4_data, fork_34_out3_data, fork_34_out2_data, fork_34_out1_data}), .valid_out_bus({fork_34_out6_valid, fork_34_out5_valid, fork_34_out4_valid, fork_34_out3_valid, fork_34_out2_valid, fork_34_out1_valid}), .ready_out_bus({fork_34_out6_ready, fork_34_out5_ready, fork_34_out4_ready, fork_34_out3_ready, fork_34_out2_ready, fork_34_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_25 (.clk(branch_25_clk), .rst(branch_25_rst), .data_in_bus({{31'b0, branch_25_in2_data}, branch_25_in1_data}), .valid_in_bus({branch_25_in2_valid, branch_25_in1_valid}), .ready_in_bus({branch_25_in2_ready, branch_25_in1_ready}), .data_out_bus({branch_25_out2_data, branch_25_out1_data}), .valid_out_bus({branch_25_out2_valid, branch_25_out1_valid}), .ready_out_bus({branch_25_out2_ready, branch_25_out1_ready}));
mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_store_op_store_1 (.clk(store_1_clk), .rst(store_1_rst), .data_in_bus({store_1_in1_data}), .address_in_bus({store_1_in2_data}), .valid_in_bus({store_1_in2_valid, store_1_in1_valid}), .ready_in_bus({store_1_in2_ready, store_1_in1_ready}), .data_out_bus({store_1_out1_data}), .address_out_bus({store_1_out2_data}), .valid_out_bus({store_1_out2_valid, store_1_out1_valid}), .ready_out_bus({store_1_out2_ready, store_1_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_41 (.clk(phiC_41_clk), .rst(phiC_41_rst), .data_in_bus({phiC_41_in1_data}), .valid_in_bus({phiC_41_in1_valid}), .ready_in_bus({phiC_41_in1_ready}), .data_out_bus({phiC_41_out1_data}), .valid_out_bus({phiC_41_out1_valid}), .ready_out_bus({phiC_41_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_29 (.clk(branch_29_clk), .rst(branch_29_rst), .data_in_bus({{31'b0, branch_29_in2_data}, branch_29_in1_data}), .valid_in_bus({branch_29_in2_valid, branch_29_in1_valid}), .ready_in_bus({branch_29_in2_ready, branch_29_in1_ready}), .data_out_bus({branch_29_out2_data, branch_29_out1_data}), .valid_out_bus({branch_29_out2_valid, branch_29_out1_valid}), .ready_out_bus({branch_29_out2_ready, branch_29_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_22 (.clk(branch_22_clk), .rst(branch_22_rst), .data_in_bus({{31'b0, branch_22_in2_data}, branch_22_in1_data}), .valid_in_bus({branch_22_in2_valid, branch_22_in1_valid}), .ready_in_bus({branch_22_in2_ready, branch_22_in1_ready}), .data_out_bus({branch_22_out2_data, branch_22_out1_data}), .valid_out_bus({branch_22_out2_valid, branch_22_out1_valid}), .ready_out_bus({branch_22_out2_ready, branch_22_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_1 (.clk(fork_1_clk), .rst(fork_1_rst), .data_in_bus({fork_1_in1_data}), .valid_in_bus({fork_1_in1_valid}), .ready_in_bus({fork_1_in1_ready}), .data_out_bus({fork_1_out2_data, fork_1_out1_data}), .valid_out_bus({fork_1_out2_valid, fork_1_out1_valid}), .ready_out_bus({fork_1_out2_ready, fork_1_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(12), .DATA_SIZE(32)) mc_load_op_load_47 (.clk(load_47_clk), .rst(load_47_rst), .data_in_bus({load_47_in1_data}), .address_in_bus({load_47_in2_data}), .valid_in_bus({load_47_in2_valid, load_47_in1_valid}), .ready_in_bus({load_47_in2_ready, load_47_in1_ready}), .data_out_bus({load_47_out1_data}), .address_out_bus({load_47_out2_data}), .valid_out_bus({load_47_out2_valid, load_47_out1_valid}), .ready_out_bus({load_47_out2_ready, load_47_out1_ready}));
shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(11), .DATA_OUT_SIZE(11)) shl_op_shl_84 (.clk(shl_84_clk), .rst(shl_84_rst), .data_in_bus({shl_84_in2_data, shl_84_in1_data}), .valid_in_bus({shl_84_in2_valid, shl_84_in1_valid}), .ready_in_bus({shl_84_in2_ready, shl_84_in1_ready}), .data_out_bus({shl_84_out1_data}), .valid_out_bus({shl_84_out1_valid}), .ready_out_bus({shl_84_out1_ready}));
mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_63 (.clk(phi_63_clk), .rst(phi_63_rst), .data_in_bus({{5'b0, phi_63_in1_data}, phi_63_in3_data, phi_63_in2_data}), .valid_in_bus({phi_63_in1_valid, phi_63_in3_valid, phi_63_in2_valid}), .ready_in_bus({phi_63_in1_ready, phi_63_in3_ready, phi_63_in2_ready}), .data_out_bus({phi_63_out1_data}), .valid_out_bus({phi_63_out1_valid}), .ready_out_bus({phi_63_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n23 (.clk(phi_n23_clk), .rst(phi_n23_rst), .data_in_bus({phi_n23_in1_data}), .valid_in_bus({phi_n23_in1_valid}), .ready_in_bus({phi_n23_in1_ready}), .data_out_bus({phi_n23_out1_data}), .valid_out_bus({phi_n23_out1_valid}), .ready_out_bus({phi_n23_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_40 (.clk(phiC_40_clk), .rst(phiC_40_rst), .data_in_bus({phiC_40_in1_data}), .valid_in_bus({phiC_40_in1_valid}), .ready_in_bus({phiC_40_in1_ready}), .data_out_bus({phiC_40_out1_data}), .valid_out_bus({phiC_40_out1_valid}), .ready_out_bus({phiC_40_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_15 (.clk(branch_15_clk), .rst(branch_15_rst), .data_in_bus({{31'b0, branch_15_in2_data}, branch_15_in1_data}), .valid_in_bus({branch_15_in2_valid, branch_15_in1_valid}), .ready_in_bus({branch_15_in2_ready, branch_15_in1_ready}), .data_out_bus({branch_15_out2_data, branch_15_out1_data}), .valid_out_bus({branch_15_out2_valid, branch_15_out1_valid}), .ready_out_bus({branch_15_out2_ready, branch_15_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_26 (.clk(sink_26_clk), .rst(sink_26_rst), .data_in_bus({sink_26_in1_data}), .valid_in_bus({sink_26_in1_valid}), .ready_in_bus({sink_26_in1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_24 (.clk(cst_24_clk), .rst(cst_24_rst), .data_in_bus({6'd32}), .valid_in_bus({cst_24_in1_valid}), .ready_in_bus({cst_24_in1_ready}), .data_out_bus({cst_24_out1_data}), .valid_out_bus({cst_24_out1_valid}), .ready_out_bus({cst_24_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n13 (.clk(phi_n13_clk), .rst(phi_n13_rst), .data_in_bus({phi_n13_in1_data}), .valid_in_bus({phi_n13_in1_valid}), .ready_in_bus({phi_n13_in1_ready}), .data_out_bus({phi_n13_out1_data}), .valid_out_bus({phi_n13_out1_valid}), .ready_out_bus({phi_n13_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_27 (.clk(branch_27_clk), .rst(branch_27_rst), .data_in_bus({{31'b0, branch_27_in2_data}, branch_27_in1_data}), .valid_in_bus({branch_27_in2_valid, branch_27_in1_valid}), .ready_in_bus({branch_27_in2_ready, branch_27_in1_ready}), .data_out_bus({branch_27_out2_data, branch_27_out1_data}), .valid_out_bus({branch_27_out2_valid, branch_27_out1_valid}), .ready_out_bus({branch_27_out2_ready, branch_27_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_14 (.clk(sink_14_clk), .rst(sink_14_rst), .data_in_bus({sink_14_in1_data}), .valid_in_bus({sink_14_in1_valid}), .ready_in_bus({sink_14_in1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n6 (.clk(phi_n6_clk), .rst(phi_n6_rst), .data_in_bus({phi_n6_in2_data, phi_n6_in1_data}), .valid_in_bus({phi_n6_in2_valid, phi_n6_in1_valid}), .ready_in_bus({phi_n6_in2_ready, phi_n6_in1_ready}), .data_out_bus({phi_n6_out1_data}), .valid_out_bus({phi_n6_out1_valid}), .ready_out_bus({phi_n6_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_17 (.clk(branch_17_clk), .rst(branch_17_rst), .data_in_bus({{31'b0, branch_17_in2_data}, branch_17_in1_data}), .valid_in_bus({branch_17_in2_valid, branch_17_in1_valid}), .ready_in_bus({branch_17_in2_ready, branch_17_in1_ready}), .data_out_bus({branch_17_out2_data, branch_17_out1_data}), .valid_out_bus({branch_17_out2_valid, branch_17_out1_valid}), .ready_out_bus({branch_17_out2_ready, branch_17_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_24 (.clk(sink_24_clk), .rst(sink_24_rst), .data_in_bus({sink_24_in1_data}), .valid_in_bus({sink_24_in1_valid}), .ready_in_bus({sink_24_in1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_16 (.clk(sink_16_clk), .rst(sink_16_rst), .data_in_bus({sink_16_in1_data}), .valid_in_bus({sink_16_in1_valid}), .ready_in_bus({sink_16_in1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_53 (.clk(forkC_53_clk), .rst(forkC_53_rst), .data_in_bus({forkC_53_in1_data}), .valid_in_bus({forkC_53_in1_valid}), .ready_in_bus({forkC_53_in1_ready}), .data_out_bus({forkC_53_out2_data, forkC_53_out1_data}), .valid_out_bus({forkC_53_out2_valid, forkC_53_out1_valid}), .ready_out_bus({forkC_53_out2_ready, forkC_53_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_41 (.clk(fork_41_clk), .rst(fork_41_rst), .data_in_bus({fork_41_in1_data}), .valid_in_bus({fork_41_in1_valid}), .ready_in_bus({fork_41_in1_ready}), .data_out_bus({fork_41_out5_data, fork_41_out4_data, fork_41_out3_data, fork_41_out2_data, fork_41_out1_data}), .valid_out_bus({fork_41_out5_valid, fork_41_out4_valid, fork_41_out3_valid, fork_41_out2_valid, fork_41_out1_valid}), .ready_out_bus({fork_41_out5_ready, fork_41_out4_ready, fork_41_out3_ready, fork_41_out2_ready, fork_41_out1_ready}));
cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_36 (.clk(phiC_36_clk), .rst(phiC_36_rst), .data_in_bus({phiC_36_in2_data, phiC_36_in1_data}), .valid_in_bus({phiC_36_in2_valid, phiC_36_in1_valid}), .ready_in_bus({phiC_36_in2_ready, phiC_36_in1_ready}), .data_out_bus({phiC_36_out2_data, phiC_36_out1_data}), .valid_out_bus({phiC_36_out2_valid, phiC_36_out1_valid}), .ready_out_bus({phiC_36_out2_ready, phiC_36_out1_ready}));
mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_store_op_store_3 (.clk(store_3_clk), .rst(store_3_rst), .data_in_bus({store_3_in1_data}), .address_in_bus({store_3_in2_data}), .valid_in_bus({store_3_in2_valid, store_3_in1_valid}), .ready_in_bus({store_3_in2_ready, store_3_in1_ready}), .data_out_bus({store_3_out1_data}), .address_out_bus({store_3_out2_data}), .valid_out_bus({store_3_out2_valid, store_3_out1_valid}), .ready_out_bus({store_3_out2_ready, store_3_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_5 (.clk(sink_5_clk), .rst(sink_5_rst), .data_in_bus({sink_5_in1_data}), .valid_in_bus({sink_5_in1_valid}), .ready_in_bus({sink_5_in1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_0 (.clk(sink_0_clk), .rst(sink_0_rst), .data_in_bus({sink_0_in1_data}), .valid_in_bus({sink_0_in1_valid}), .ready_in_bus({sink_0_in1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block2 (.clk(brCst_block2_clk), .rst(brCst_block2_rst), .data_in_bus({1'd1}), .valid_in_bus({brCst_block2_in1_valid}), .ready_in_bus({brCst_block2_in1_ready}), .data_out_bus({brCst_block2_out1_data}), .valid_out_bus({brCst_block2_out1_valid}), .ready_out_bus({brCst_block2_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_18 (.clk(branch_18_clk), .rst(branch_18_rst), .data_in_bus({{branch_18_in2_data}, branch_18_in1_data}), .valid_in_bus({branch_18_in2_valid, branch_18_in1_valid}), .ready_in_bus({branch_18_in2_ready, branch_18_in1_ready}), .data_out_bus({branch_18_out2_data, branch_18_out1_data}), .valid_out_bus({branch_18_out2_valid, branch_18_out1_valid}), .ready_out_bus({branch_18_out2_ready, branch_18_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_23 (.clk(branch_23_clk), .rst(branch_23_rst), .data_in_bus({{5'b0, branch_23_in2_data}, branch_23_in1_data}), .valid_in_bus({branch_23_in2_valid, branch_23_in1_valid}), .ready_in_bus({branch_23_in2_ready, branch_23_in1_ready}), .data_out_bus({branch_23_out2_data, branch_23_out1_data}), .valid_out_bus({branch_23_out2_valid, branch_23_out1_valid}), .ready_out_bus({branch_23_out2_ready, branch_23_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_6 (.clk(cst_6_clk), .rst(cst_6_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_6_in1_valid}), .ready_in_bus({cst_6_in1_ready}), .data_out_bus({cst_6_out1_data}), .valid_out_bus({cst_6_out1_valid}), .ready_out_bus({cst_6_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(12), .DATA_OUT_SIZE(12)) add_op_add_26 (.clk(add_26_clk), .rst(add_26_rst), .data_in_bus({add_26_in2_data, add_26_in1_data}), .valid_in_bus({add_26_in2_valid, add_26_in1_valid}), .ready_in_bus({add_26_in2_ready, add_26_in1_ready}), .data_out_bus({add_26_out1_data}), .valid_out_bus({add_26_out1_valid}), .ready_out_bus({add_26_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) OEHB_Buffer_16 (.clk(Buffer_16_clk), .rst(Buffer_16_rst), .data_in_bus({Buffer_16_in1_data}), .valid_in_bus({Buffer_16_in1_valid}), .ready_in_bus({Buffer_16_in1_ready}), .data_out_bus({Buffer_16_out1_data}), .valid_out_bus({Buffer_16_out1_valid}), .ready_out_bus({Buffer_16_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_35 (.clk(phiC_35_clk), .rst(phiC_35_rst), .data_in_bus({phiC_35_in1_data}), .valid_in_bus({phiC_35_in1_valid}), .ready_in_bus({phiC_35_in1_ready}), .data_out_bus({phiC_35_out1_data}), .valid_out_bus({phiC_35_out1_valid}), .ready_out_bus({phiC_35_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_40 (.clk(branch_40_clk), .rst(branch_40_rst), .data_in_bus({{31'b0, branch_40_in2_data}, branch_40_in1_data}), .valid_in_bus({branch_40_in2_valid, branch_40_in1_valid}), .ready_in_bus({branch_40_in2_ready, branch_40_in1_ready}), .data_out_bus({branch_40_out2_data, branch_40_out1_data}), .valid_out_bus({branch_40_out2_valid, branch_40_out1_valid}), .ready_out_bus({branch_40_out2_ready, branch_40_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_1 (.clk(source_1_clk), .rst(source_1_rst), .data_out_bus({source_1_out1_data}), .valid_out_bus({source_1_out1_valid}), .ready_out_bus({source_1_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_69 (.clk(load_69_clk), .rst(load_69_rst), .data_in_bus({load_69_in1_data}), .address_in_bus({load_69_in2_data}), .valid_in_bus({load_69_in2_valid, load_69_in1_valid}), .ready_in_bus({load_69_in2_ready, load_69_in1_ready}), .data_out_bus({load_69_out1_data}), .address_out_bus({load_69_out2_data}), .valid_out_bus({load_69_out2_valid, load_69_out1_valid}), .ready_out_bus({load_69_out2_ready, load_69_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_42 (.clk(branch_42_clk), .rst(branch_42_rst), .data_in_bus({{5'b0, branch_42_in2_data}, branch_42_in1_data}), .valid_in_bus({branch_42_in2_valid, branch_42_in1_valid}), .ready_in_bus({branch_42_in2_ready, branch_42_in1_ready}), .data_out_bus({branch_42_out2_data, branch_42_out1_data}), .valid_out_bus({branch_42_out2_valid, branch_42_out1_valid}), .ready_out_bus({branch_42_out2_ready, branch_42_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_19 (.clk(branch_19_clk), .rst(branch_19_rst), .data_in_bus({{31'b0, branch_19_in2_data}, branch_19_in1_data}), .valid_in_bus({branch_19_in2_valid, branch_19_in1_valid}), .ready_in_bus({branch_19_in2_ready, branch_19_in1_ready}), .data_out_bus({branch_19_out2_data, branch_19_out1_data}), .valid_out_bus({branch_19_out2_valid, branch_19_out1_valid}), .ready_out_bus({branch_19_out2_ready, branch_19_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block9 (.clk(brCst_block9_clk), .rst(brCst_block9_rst), .data_in_bus({1'd1}), .valid_in_bus({brCst_block9_in1_valid}), .ready_in_bus({brCst_block9_in1_ready}), .data_out_bus({brCst_block9_out1_data}), .valid_out_bus({brCst_block9_out1_valid}), .ready_out_bus({brCst_block9_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_23 (.clk(fork_23_clk), .rst(fork_23_rst), .data_in_bus({fork_23_in1_data}), .valid_in_bus({fork_23_in1_valid}), .ready_in_bus({fork_23_in1_ready}), .data_out_bus({fork_23_out2_data, fork_23_out1_data}), .valid_out_bus({fork_23_out2_valid, fork_23_out1_valid}), .ready_out_bus({fork_23_out2_ready, fork_23_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_26 (.clk(cst_26_clk), .rst(cst_26_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_26_in1_valid}), .ready_in_bus({cst_26_in1_ready}), .data_out_bus({cst_26_out1_data}), .valid_out_bus({cst_26_out1_valid}), .ready_out_bus({cst_26_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_55 (.clk(branchC_55_clk), .rst(branchC_55_rst), .data_in_bus({{branchC_55_in2_data}, branchC_55_in1_data}), .valid_in_bus({branchC_55_in2_valid, branchC_55_in1_valid}), .ready_in_bus({branchC_55_in2_ready, branchC_55_in1_ready}), .data_out_bus({branchC_55_out2_data, branchC_55_out1_data}), .valid_out_bus({branchC_55_out2_valid, branchC_55_out1_valid}), .ready_out_bus({branchC_55_out2_ready, branchC_55_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_51 (.clk(branchC_51_clk), .rst(branchC_51_rst), .data_in_bus({{branchC_51_in2_data}, branchC_51_in1_data}), .valid_in_bus({branchC_51_in2_valid, branchC_51_in1_valid}), .ready_in_bus({branchC_51_in2_ready, branchC_51_in1_ready}), .data_out_bus({branchC_51_out2_data, branchC_51_out1_data}), .valid_out_bus({branchC_51_out2_valid, branchC_51_out1_valid}), .ready_out_bus({branchC_51_out2_ready, branchC_51_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n12 (.clk(phi_n12_clk), .rst(phi_n12_rst), .data_in_bus({phi_n12_in1_data}), .valid_in_bus({phi_n12_in1_valid}), .ready_in_bus({phi_n12_in1_ready}), .data_out_bus({phi_n12_out1_data}), .valid_out_bus({phi_n12_out1_valid}), .ready_out_bus({phi_n12_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_12 (.clk(branch_12_clk), .rst(branch_12_rst), .data_in_bus({{31'b0, branch_12_in2_data}, branch_12_in1_data}), .valid_in_bus({branch_12_in2_valid, branch_12_in1_valid}), .ready_in_bus({branch_12_in2_ready, branch_12_in1_ready}), .data_out_bus({branch_12_out2_data, branch_12_out1_data}), .valid_out_bus({branch_12_out2_valid, branch_12_out1_valid}), .ready_out_bus({branch_12_out2_ready, branch_12_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(12), .DATA_OUT_SIZE(12)) add_op_add_5 (.clk(add_5_clk), .rst(add_5_rst), .data_in_bus({add_5_in2_data, add_5_in1_data}), .valid_in_bus({add_5_in2_valid, add_5_in1_valid}), .ready_in_bus({add_5_in2_ready, add_5_in1_ready}), .data_out_bus({add_5_out1_data}), .valid_out_bus({add_5_out1_valid}), .ready_out_bus({add_5_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_10 (.clk(branch_10_clk), .rst(branch_10_rst), .data_in_bus({{31'b0, branch_10_in2_data}, branch_10_in1_data}), .valid_in_bus({branch_10_in2_valid, branch_10_in1_valid}), .ready_in_bus({branch_10_in2_ready, branch_10_in1_ready}), .data_out_bus({branch_10_out2_data, branch_10_out1_data}), .valid_out_bus({branch_10_out2_valid, branch_10_out1_valid}), .ready_out_bus({branch_10_out2_ready, branch_10_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_0 (.clk(source_0_clk), .rst(source_0_rst), .data_out_bus({source_0_out1_data}), .valid_out_bus({source_0_out1_valid}), .ready_out_bus({source_0_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_31 (.clk(branch_31_clk), .rst(branch_31_rst), .data_in_bus({{31'b0, branch_31_in2_data}, branch_31_in1_data}), .valid_in_bus({branch_31_in2_valid, branch_31_in1_valid}), .ready_in_bus({branch_31_in2_ready, branch_31_in1_ready}), .data_out_bus({branch_31_out2_data, branch_31_out1_data}), .valid_out_bus({branch_31_out2_valid, branch_31_out1_valid}), .ready_out_bus({branch_31_out2_ready, branch_31_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_19 (.clk(cst_19_clk), .rst(cst_19_rst), .data_in_bus({1'd0}), .valid_in_bus({cst_19_in1_valid}), .ready_in_bus({cst_19_in1_ready}), .data_out_bus({cst_19_out1_data}), .valid_out_bus({cst_19_out1_valid}), .ready_out_bus({cst_19_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n9 (.clk(phi_n9_clk), .rst(phi_n9_rst), .data_in_bus({phi_n9_in1_data}), .valid_in_bus({phi_n9_in1_valid}), .ready_in_bus({phi_n9_in1_ready}), .data_out_bus({phi_n9_out1_data}), .valid_out_bus({phi_n9_out1_valid}), .ready_out_bus({phi_n9_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_46 (.clk(branchC_46_clk), .rst(branchC_46_rst), .data_in_bus({{branchC_46_in2_data}, branchC_46_in1_data}), .valid_in_bus({branchC_46_in2_valid, branchC_46_in1_valid}), .ready_in_bus({branchC_46_in2_ready, branchC_46_in1_ready}), .data_out_bus({branchC_46_out2_data, branchC_46_out1_data}), .valid_out_bus({branchC_46_out2_valid, branchC_46_out1_valid}), .ready_out_bus({branchC_46_out2_ready, branchC_46_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_36 (.clk(fork_36_clk), .rst(fork_36_rst), .data_in_bus({fork_36_in1_data}), .valid_in_bus({fork_36_in1_valid}), .ready_in_bus({fork_36_in1_ready}), .data_out_bus({fork_36_out4_data, fork_36_out3_data, fork_36_out2_data, fork_36_out1_data}), .valid_out_bus({fork_36_out4_valid, fork_36_out3_valid, fork_36_out2_valid, fork_36_out1_valid}), .ready_out_bus({fork_36_out4_ready, fork_36_out3_ready, fork_36_out2_ready, fork_36_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_5 (.clk(cst_5_clk), .rst(cst_5_rst), .data_in_bus({6'd32}), .valid_in_bus({cst_5_in1_valid}), .ready_in_bus({cst_5_in1_ready}), .data_out_bus({cst_5_out1_data}), .valid_out_bus({cst_5_out1_valid}), .ready_out_bus({cst_5_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n24 (.clk(phi_n24_clk), .rst(phi_n24_rst), .data_in_bus({phi_n24_in1_data}), .valid_in_bus({phi_n24_in1_valid}), .ready_in_bus({phi_n24_in1_ready}), .data_out_bus({phi_n24_out1_data}), .valid_out_bus({phi_n24_out1_valid}), .ready_out_bus({phi_n24_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_5 (.clk(Buffer_5_clk), .rst(Buffer_5_rst), .data_in_bus({Buffer_5_in1_data}), .valid_in_bus({Buffer_5_in1_valid}), .ready_in_bus({Buffer_5_in1_ready}), .data_out_bus({Buffer_5_out1_data}), .valid_out_bus({Buffer_5_out1_valid}), .ready_out_bus({Buffer_5_out1_ready}));
mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_41 (.clk(phi_41_clk), .rst(phi_41_rst), .data_in_bus({{31'b0, phi_41_in1_data}, phi_41_in3_data, phi_41_in2_data}), .valid_in_bus({phi_41_in1_valid, phi_41_in3_valid, phi_41_in2_valid}), .ready_in_bus({phi_41_in1_ready, phi_41_in3_ready, phi_41_in2_ready}), .data_out_bus({phi_41_out1_data}), .valid_out_bus({phi_41_out1_valid}), .ready_out_bus({phi_41_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n8 (.clk(phi_n8_clk), .rst(phi_n8_rst), .data_in_bus({phi_n8_in1_data}), .valid_in_bus({phi_n8_in1_valid}), .ready_in_bus({phi_n8_in1_ready}), .data_out_bus({phi_n8_out1_data}), .valid_out_bus({phi_n8_out1_valid}), .ready_out_bus({phi_n8_out1_ready}));
cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_39 (.clk(phiC_39_clk), .rst(phiC_39_rst), .data_in_bus({phiC_39_in2_data, phiC_39_in1_data}), .valid_in_bus({phiC_39_in2_valid, phiC_39_in1_valid}), .ready_in_bus({phiC_39_in2_ready, phiC_39_in1_ready}), .data_out_bus({phiC_39_out2_data, phiC_39_out1_data}), .valid_out_bus({phiC_39_out2_valid, phiC_39_out1_valid}), .ready_out_bus({phiC_39_out2_ready, phiC_39_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_27 (.clk(sink_27_clk), .rst(sink_27_rst), .data_in_bus({sink_27_in1_data}), .valid_in_bus({sink_27_in1_valid}), .ready_in_bus({sink_27_in1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_22 (.clk(fork_22_clk), .rst(fork_22_rst), .data_in_bus({fork_22_in1_data}), .valid_in_bus({fork_22_in1_valid}), .ready_in_bus({fork_22_in1_ready}), .data_out_bus({fork_22_out2_data, fork_22_out1_data}), .valid_out_bus({fork_22_out2_valid, fork_22_out1_valid}), .ready_out_bus({fork_22_out2_ready, fork_22_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_31 (.clk(phiC_31_clk), .rst(phiC_31_rst), .data_in_bus({phiC_31_in1_data}), .valid_in_bus({phiC_31_in1_valid}), .ready_in_bus({phiC_31_in1_ready}), .data_out_bus({phiC_31_out1_data}), .valid_out_bus({phiC_31_out1_valid}), .ready_out_bus({phiC_31_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_6 (.clk(sink_6_clk), .rst(sink_6_rst), .data_in_bus({sink_6_in1_data}), .valid_in_bus({sink_6_in1_valid}), .ready_in_bus({sink_6_in1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_10 (.clk(sink_10_clk), .rst(sink_10_rst), .data_in_bus({sink_10_in1_data}), .valid_in_bus({sink_10_in1_valid}), .ready_in_bus({sink_10_in1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_54 (.clk(forkC_54_clk), .rst(forkC_54_rst), .data_in_bus({forkC_54_in1_data}), .valid_in_bus({forkC_54_in1_valid}), .ready_in_bus({forkC_54_in1_ready}), .data_out_bus({forkC_54_out3_data, forkC_54_out2_data, forkC_54_out1_data}), .valid_out_bus({forkC_54_out3_valid, forkC_54_out2_valid, forkC_54_out1_valid}), .ready_out_bus({forkC_54_out3_ready, forkC_54_out2_ready, forkC_54_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_31 (.clk(fork_31_clk), .rst(fork_31_rst), .data_in_bus({fork_31_in1_data}), .valid_in_bus({fork_31_in1_valid}), .ready_in_bus({fork_31_in1_ready}), .data_out_bus({fork_31_out5_data, fork_31_out4_data, fork_31_out3_data, fork_31_out2_data, fork_31_out1_data}), .valid_out_bus({fork_31_out5_valid, fork_31_out4_valid, fork_31_out3_valid, fork_31_out2_valid, fork_31_out1_valid}), .ready_out_bus({fork_31_out5_ready, fork_31_out4_ready, fork_31_out3_ready, fork_31_out2_ready, fork_31_out1_ready}));
mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_1 (.clk(phi_1_clk), .rst(phi_1_rst), .data_in_bus({{5'b0, phi_1_in1_data}, phi_1_in3_data, phi_1_in2_data}), .valid_in_bus({phi_1_in1_valid, phi_1_in3_valid, phi_1_in2_valid}), .ready_in_bus({phi_1_in1_ready, phi_1_in3_ready, phi_1_in2_ready}), .data_out_bus({phi_1_out1_data}), .valid_out_bus({phi_1_out1_valid}), .ready_out_bus({phi_1_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(12), .DATA_OUT_SIZE(12)) add_op_add_85 (.clk(add_85_clk), .rst(add_85_rst), .data_in_bus({add_85_in2_data, add_85_in1_data}), .valid_in_bus({add_85_in2_valid, add_85_in1_valid}), .ready_in_bus({add_85_in2_ready, add_85_in1_ready}), .data_out_bus({add_85_out1_data}), .valid_out_bus({add_85_out1_valid}), .ready_out_bus({add_85_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_27 (.clk(fork_27_clk), .rst(fork_27_rst), .data_in_bus({fork_27_in1_data}), .valid_in_bus({fork_27_in1_valid}), .ready_in_bus({fork_27_in1_ready}), .data_out_bus({fork_27_out2_data, fork_27_out1_data}), .valid_out_bus({fork_27_out2_valid, fork_27_out1_valid}), .ready_out_bus({fork_27_out2_ready, fork_27_out1_ready}));
cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_32 (.clk(phiC_32_clk), .rst(phiC_32_rst), .data_in_bus({phiC_32_in2_data, phiC_32_in1_data}), .valid_in_bus({phiC_32_in2_valid, phiC_32_in1_valid}), .ready_in_bus({phiC_32_in2_ready, phiC_32_in1_ready}), .data_out_bus({phiC_32_out2_data, phiC_32_out1_data}), .valid_out_bus({phiC_32_out2_valid, phiC_32_out1_valid}), .ready_out_bus({phiC_32_out2_ready, phiC_32_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block11 (.clk(brCst_block11_clk), .rst(brCst_block11_rst), .data_in_bus({1'd1}), .valid_in_bus({brCst_block11_in1_valid}), .ready_in_bus({brCst_block11_in1_ready}), .data_out_bus({brCst_block11_out1_data}), .valid_out_bus({brCst_block11_out1_valid}), .ready_out_bus({brCst_block11_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_11 (.clk(source_11_clk), .rst(source_11_rst), .data_out_bus({source_11_out1_data}), .valid_out_bus({source_11_out1_valid}), .ready_out_bus({source_11_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_7 (.clk(sink_7_clk), .rst(sink_7_rst), .data_in_bus({sink_7_in1_data}), .valid_in_bus({sink_7_in1_valid}), .ready_in_bus({sink_7_in1_ready}));
mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(16), .DATA_OUT_SIZE(32)) mul_op_mul_48 (.clk(mul_48_clk), .rst(mul_48_rst), .data_in_bus({mul_48_in2_data, mul_48_in1_data}), .valid_in_bus({mul_48_in2_valid, mul_48_in1_valid}), .ready_in_bus({mul_48_in2_ready, mul_48_in1_ready}), .data_out_bus({mul_48_out1_data}), .valid_out_bus({mul_48_out1_valid}), .ready_out_bus({mul_48_out1_ready}));
cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_38 (.clk(phiC_38_clk), .rst(phiC_38_rst), .data_in_bus({phiC_38_in2_data, phiC_38_in1_data}), .valid_in_bus({phiC_38_in2_valid, phiC_38_in1_valid}), .ready_in_bus({phiC_38_in2_ready, phiC_38_in1_ready}), .data_out_bus({phiC_38_out2_data, phiC_38_out1_data}), .valid_out_bus({phiC_38_out2_valid, phiC_38_out1_valid}), .ready_out_bus({phiC_38_out2_ready, phiC_38_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_8 (.clk(sink_8_clk), .rst(sink_8_rst), .data_in_bus({sink_8_in1_data}), .valid_in_bus({sink_8_in1_valid}), .ready_in_bus({sink_8_in1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_21 (.clk(cst_21_clk), .rst(cst_21_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_21_in1_valid}), .ready_in_bus({cst_21_in1_ready}), .data_out_bus({cst_21_out1_data}), .valid_out_bus({cst_21_out1_valid}), .ready_out_bus({cst_21_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_54 (.clk(branchC_54_clk), .rst(branchC_54_rst), .data_in_bus({{branchC_54_in2_data}, branchC_54_in1_data}), .valid_in_bus({branchC_54_in2_valid, branchC_54_in1_valid}), .ready_in_bus({branchC_54_in2_ready, branchC_54_in1_ready}), .data_out_bus({branchC_54_out2_data, branchC_54_out1_data}), .valid_out_bus({branchC_54_out2_valid, branchC_54_out1_valid}), .ready_out_bus({branchC_54_out2_ready, branchC_54_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_9 (.clk(branch_9_clk), .rst(branch_9_rst), .data_in_bus({{31'b0, branch_9_in2_data}, branch_9_in1_data}), .valid_in_bus({branch_9_in2_valid, branch_9_in1_valid}), .ready_in_bus({branch_9_in2_ready, branch_9_in1_ready}), .data_out_bus({branch_9_out2_data, branch_9_out1_data}), .valid_out_bus({branch_9_out2_valid, branch_9_out1_valid}), .ready_out_bus({branch_9_out2_ready, branch_9_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n3 (.clk(phi_n3_clk), .rst(phi_n3_rst), .data_in_bus({phi_n3_in1_data}), .valid_in_bus({phi_n3_in1_valid}), .ready_in_bus({phi_n3_in1_ready}), .data_out_bus({phi_n3_out1_data}), .valid_out_bus({phi_n3_out1_valid}), .ready_out_bus({phi_n3_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_16 (.clk(branch_16_clk), .rst(branch_16_rst), .data_in_bus({{31'b0, branch_16_in2_data}, branch_16_in1_data}), .valid_in_bus({branch_16_in2_valid, branch_16_in1_valid}), .ready_in_bus({branch_16_in2_ready, branch_16_in1_ready}), .data_out_bus({branch_16_out2_data, branch_16_out1_data}), .valid_out_bus({branch_16_out2_valid, branch_16_out1_valid}), .ready_out_bus({branch_16_out2_ready, branch_16_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n25 (.clk(phi_n25_clk), .rst(phi_n25_rst), .data_in_bus({phi_n25_in1_data}), .valid_in_bus({phi_n25_in1_valid}), .ready_in_bus({phi_n25_in1_ready}), .data_out_bus({phi_n25_out1_data}), .valid_out_bus({phi_n25_out1_valid}), .ready_out_bus({phi_n25_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_45 (.clk(branch_45_clk), .rst(branch_45_rst), .data_in_bus({{5'b0, branch_45_in2_data}, branch_45_in1_data}), .valid_in_bus({branch_45_in2_valid, branch_45_in1_valid}), .ready_in_bus({branch_45_in2_ready, branch_45_in1_ready}), .data_out_bus({branch_45_out2_data, branch_45_out1_data}), .valid_out_bus({branch_45_out2_valid, branch_45_out1_valid}), .ready_out_bus({branch_45_out2_ready, branch_45_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n21 (.clk(phi_n21_clk), .rst(phi_n21_rst), .data_in_bus({phi_n21_in1_data}), .valid_in_bus({phi_n21_in1_valid}), .ready_in_bus({phi_n21_in1_ready}), .data_out_bus({phi_n21_out1_data}), .valid_out_bus({phi_n21_out1_valid}), .ready_out_bus({phi_n21_out1_ready}));
MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_u2 (.clk(MC_u2_clk), .rst(MC_u2_rst), .io_storeDataOut(u2_dout0), .io_storeAddrOut(u2_address0), .io_storeEnable(u2_we0), .io_loadDataIn(u2_din1), .io_loadAddrOut(u2_address1), .io_loadEnable(u2_ce1), .io_bbpValids({MC_u2_in2_valid}), .io_bb_stCountArray({MC_u2_in2_data}), .io_bbReadyToPrevs({MC_u2_in2_ready}), .io_rdPortsPrev_ready({MC_u2_in1_ready}), .io_rdPortsPrev_valid({MC_u2_in1_valid}), .io_rdPortsPrev_bits({MC_u2_in1_data}), .io_wrAddrPorts_ready({MC_u2_in3_ready}), .io_wrAddrPorts_valid({MC_u2_in3_valid}), .io_wrAddrPorts_bits({MC_u2_in3_data}), .io_wrDataPorts_ready({MC_u2_in4_ready}), .io_wrDataPorts_valid({MC_u2_in4_valid}), .io_wrDataPorts_bits({MC_u2_in4_data}), .io_rdPortsNext_ready({MC_u2_out1_ready}), .io_rdPortsNext_valid({MC_u2_out1_valid}), .io_rdPortsNext_bits({MC_u2_out1_data}), .io_Empty_Valid({MC_u2_out2_valid}), .io_Empty_Ready({MC_u2_out2_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) OEHB_Buffer_27 (.clk(Buffer_27_clk), .rst(Buffer_27_rst), .data_in_bus({Buffer_27_in1_data}), .valid_in_bus({Buffer_27_in1_valid}), .ready_in_bus({Buffer_27_in1_ready}), .data_out_bus({Buffer_27_out1_data}), .valid_out_bus({Buffer_27_out1_valid}), .ready_out_bus({Buffer_27_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_70 (.clk(add_70_clk), .rst(add_70_rst), .data_in_bus({add_70_in2_data, add_70_in1_data}), .valid_in_bus({add_70_in2_valid, add_70_in1_valid}), .ready_in_bus({add_70_in2_ready, add_70_in1_ready}), .data_out_bus({add_70_out1_data}), .valid_out_bus({add_70_out1_valid}), .ready_out_bus({add_70_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_18 (.clk(sink_18_clk), .rst(sink_18_rst), .data_in_bus({sink_18_in1_data}), .valid_in_bus({sink_18_in1_valid}), .ready_in_bus({sink_18_in1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) OEHB_Buffer_10 (.clk(Buffer_10_clk), .rst(Buffer_10_rst), .data_in_bus({Buffer_10_in1_data}), .valid_in_bus({Buffer_10_in1_valid}), .ready_in_bus({Buffer_10_in1_ready}), .data_out_bus({Buffer_10_out1_data}), .valid_out_bus({Buffer_10_out1_valid}), .ready_out_bus({Buffer_10_out1_ready}));
icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_33 (.clk(icmp_33_clk), .rst(icmp_33_rst), .data_in_bus({icmp_33_in2_data, icmp_33_in1_data}), .valid_in_bus({icmp_33_in2_valid, icmp_33_in1_valid}), .ready_in_bus({icmp_33_in2_ready, icmp_33_in1_ready}), .data_out_bus({icmp_33_out1_data}), .valid_out_bus({icmp_33_out1_valid}), .ready_out_bus({icmp_33_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_12 (.clk(Buffer_12_clk), .rst(Buffer_12_rst), .data_in_bus({Buffer_12_in1_data}), .valid_in_bus({Buffer_12_in1_valid}), .ready_in_bus({Buffer_12_in1_ready}), .data_out_bus({Buffer_12_out1_data}), .valid_out_bus({Buffer_12_out1_valid}), .ready_out_bus({Buffer_12_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_95 (.clk(add_95_clk), .rst(add_95_rst), .data_in_bus({add_95_in2_data, add_95_in1_data}), .valid_in_bus({add_95_in2_valid, add_95_in1_valid}), .ready_in_bus({add_95_in2_ready, add_95_in1_ready}), .data_out_bus({add_95_out1_data}), .valid_out_bus({add_95_out1_valid}), .ready_out_bus({add_95_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_23 (.clk(cst_23_clk), .rst(cst_23_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_23_in1_valid}), .ready_in_bus({cst_23_in1_ready}), .data_out_bus({cst_23_out1_data}), .valid_out_bus({cst_23_out1_valid}), .ready_out_bus({cst_23_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_11 (.clk(branch_11_clk), .rst(branch_11_rst), .data_in_bus({{5'b0, branch_11_in2_data}, branch_11_in1_data}), .valid_in_bus({branch_11_in2_valid, branch_11_in1_valid}), .ready_in_bus({branch_11_in2_ready, branch_11_in1_ready}), .data_out_bus({branch_11_out2_data, branch_11_out1_data}), .valid_out_bus({branch_11_out2_valid, branch_11_out1_valid}), .ready_out_bus({branch_11_out2_ready, branch_11_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_50 (.clk(branchC_50_clk), .rst(branchC_50_rst), .data_in_bus({{branchC_50_in2_data}, branchC_50_in1_data}), .valid_in_bus({branchC_50_in2_valid, branchC_50_in1_valid}), .ready_in_bus({branchC_50_in2_ready, branchC_50_in1_ready}), .data_out_bus({branchC_50_out2_data, branchC_50_out1_data}), .valid_out_bus({branchC_50_out2_valid, branchC_50_out1_valid}), .ready_out_bus({branchC_50_out2_ready, branchC_50_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_8 (.clk(cst_8_clk), .rst(cst_8_rst), .data_in_bus({1'd0}), .valid_in_bus({cst_8_in1_valid}), .ready_in_bus({cst_8_in1_ready}), .data_out_bus({cst_8_out1_data}), .valid_out_bus({cst_8_out1_valid}), .ready_out_bus({cst_8_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_44 (.clk(forkC_44_clk), .rst(forkC_44_rst), .data_in_bus({forkC_44_in1_data}), .valid_in_bus({forkC_44_in1_valid}), .ready_in_bus({forkC_44_in1_ready}), .data_out_bus({forkC_44_out3_data, forkC_44_out2_data, forkC_44_out1_data}), .valid_out_bus({forkC_44_out3_valid, forkC_44_out2_valid, forkC_44_out1_valid}), .ready_out_bus({forkC_44_out3_ready, forkC_44_out2_ready, forkC_44_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) OEHB_Buffer_7 (.clk(Buffer_7_clk), .rst(Buffer_7_rst), .data_in_bus({Buffer_7_in1_data}), .valid_in_bus({Buffer_7_in1_valid}), .ready_in_bus({Buffer_7_in1_ready}), .data_out_bus({Buffer_7_out1_data}), .valid_out_bus({Buffer_7_out1_valid}), .ready_out_bus({Buffer_7_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n27 (.clk(phi_n27_clk), .rst(phi_n27_rst), .data_in_bus({phi_n27_in2_data, phi_n27_in1_data}), .valid_in_bus({phi_n27_in2_valid, phi_n27_in1_valid}), .ready_in_bus({phi_n27_in2_ready, phi_n27_in1_ready}), .data_out_bus({phi_n27_out1_data}), .valid_out_bus({phi_n27_out1_valid}), .ready_out_bus({phi_n27_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_2 (.clk(source_2_clk), .rst(source_2_rst), .data_out_bus({source_2_out1_data}), .valid_out_bus({source_2_out1_valid}), .ready_out_bus({source_2_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_34 (.clk(branch_34_clk), .rst(branch_34_rst), .data_in_bus({{branch_34_in2_data}, branch_34_in1_data}), .valid_in_bus({branch_34_in2_valid, branch_34_in1_valid}), .ready_in_bus({branch_34_in2_ready, branch_34_in1_ready}), .data_out_bus({branch_34_out2_data, branch_34_out1_data}), .valid_out_bus({branch_34_out2_valid, branch_34_out1_valid}), .ready_out_bus({branch_34_out2_ready, branch_34_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_30 (.clk(phiC_30_clk), .rst(phiC_30_rst), .data_in_bus({phiC_30_in1_data}), .valid_in_bus({phiC_30_in1_valid}), .ready_in_bus({phiC_30_in1_ready}), .data_out_bus({phiC_30_out1_data}), .valid_out_bus({phiC_30_out1_valid}), .ready_out_bus({phiC_30_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_52 (.clk(branchC_52_clk), .rst(branchC_52_rst), .data_in_bus({{branchC_52_in2_data}, branchC_52_in1_data}), .valid_in_bus({branchC_52_in2_valid, branchC_52_in1_valid}), .ready_in_bus({branchC_52_in2_ready, branchC_52_in1_ready}), .data_out_bus({branchC_52_out2_data, branchC_52_out1_data}), .valid_out_bus({branchC_52_out2_valid, branchC_52_out1_valid}), .ready_out_bus({branchC_52_out2_ready, branchC_52_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_13 (.clk(source_13_clk), .rst(source_13_rst), .data_out_bus({source_13_out1_data}), .valid_out_bus({source_13_out1_valid}), .ready_out_bus({source_13_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_15 (.clk(cst_15_clk), .rst(cst_15_rst), .data_in_bus({1'd0}), .valid_in_bus({cst_15_in1_valid}), .ready_in_bus({cst_15_in1_ready}), .data_out_bus({cst_15_out1_data}), .valid_out_bus({cst_15_out1_valid}), .ready_out_bus({cst_15_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_59 (.clk(add_59_clk), .rst(add_59_rst), .data_in_bus({add_59_in2_data, add_59_in1_data}), .valid_in_bus({add_59_in2_valid, add_59_in1_valid}), .ready_in_bus({add_59_in2_ready, add_59_in1_ready}), .data_out_bus({add_59_out1_data}), .valid_out_bus({add_59_out1_valid}), .ready_out_bus({add_59_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_3 (.clk(branch_3_clk), .rst(branch_3_rst), .data_in_bus({{branch_3_in2_data}, branch_3_in1_data}), .valid_in_bus({branch_3_in2_valid, branch_3_in1_valid}), .ready_in_bus({branch_3_in2_ready, branch_3_in1_ready}), .data_out_bus({branch_3_out2_data, branch_3_out1_data}), .valid_out_bus({branch_3_out2_valid, branch_3_out1_valid}), .ready_out_bus({branch_3_out2_ready, branch_3_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_11 (.clk(cst_11_clk), .rst(cst_11_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_11_in1_valid}), .ready_in_bus({cst_11_in1_ready}), .data_out_bus({cst_11_out1_data}), .valid_out_bus({cst_11_out1_valid}), .ready_out_bus({cst_11_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_29 (.clk(sink_29_clk), .rst(sink_29_rst), .data_in_bus({sink_29_in1_data}), .valid_in_bus({sink_29_in1_valid}), .ready_in_bus({sink_29_in1_ready}));
mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(12), .DATA_SIZE(32)) mc_store_op_store_0 (.clk(store_0_clk), .rst(store_0_rst), .data_in_bus({store_0_in1_data}), .address_in_bus({store_0_in2_data}), .valid_in_bus({store_0_in2_valid, store_0_in1_valid}), .ready_in_bus({store_0_in2_ready, store_0_in1_ready}), .data_out_bus({store_0_out1_data}), .address_out_bus({store_0_out2_data}), .valid_out_bus({store_0_out2_valid, store_0_out1_valid}), .ready_out_bus({store_0_out2_ready, store_0_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block5 (.clk(brCst_block5_clk), .rst(brCst_block5_rst), .data_in_bus({1'd1}), .valid_in_bus({brCst_block5_in1_valid}), .ready_in_bus({brCst_block5_in1_ready}), .data_out_bus({brCst_block5_out1_data}), .valid_out_bus({brCst_block5_out1_valid}), .ready_out_bus({brCst_block5_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_14 (.clk(fork_14_clk), .rst(fork_14_rst), .data_in_bus({fork_14_in1_data}), .valid_in_bus({fork_14_in1_valid}), .ready_in_bus({fork_14_in1_ready}), .data_out_bus({fork_14_out2_data, fork_14_out1_data}), .valid_out_bus({fork_14_out2_valid, fork_14_out1_valid}), .ready_out_bus({fork_14_out2_ready, fork_14_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_2 (.clk(branch_2_clk), .rst(branch_2_rst), .data_in_bus({{31'b0, branch_2_in2_data}, branch_2_in1_data}), .valid_in_bus({branch_2_in2_valid, branch_2_in1_valid}), .ready_in_bus({branch_2_in2_ready, branch_2_in1_ready}), .data_out_bus({branch_2_out2_data, branch_2_out1_data}), .valid_out_bus({branch_2_out2_valid, branch_2_out1_valid}), .ready_out_bus({branch_2_out2_ready, branch_2_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_17 (.clk(sink_17_clk), .rst(sink_17_rst), .data_in_bus({sink_17_in1_data}), .valid_in_bus({sink_17_in1_valid}), .ready_in_bus({sink_17_in1_ready}));
endmodule
