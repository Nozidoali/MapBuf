module insertion_sort(
	input branch_8__phi_n2__valid__0__anchor__in,
	input forkC_23__brCst_block2__ready__0__anchor__in,
	input [31 : 0] fork_8__add_17__data__0__anchor__in,
	input fork_15__branch_6__valid__0__anchor__in,
	input forkC_27__branchC_26__ready__0__anchor__in,
	input [31 : 0] Buffer_55__phi_n6__data__0__anchor__in,
	input [31 : 0] fork_8__store_0__data__0__anchor__in,
	input branch_3__phi_n6__ready__0__anchor__in,
	input forkC_28__cst_8__ready__0__anchor__in,
	input forkC_23__branchC_22__ready__0__anchor__in,
	input branch_1__phi_3__ready__0__anchor__in,
	input phi_n10__branch_16__ready__0__anchor__in,
	input fork_18__branch_16__valid__0__anchor__in,
	input [31 : 0] phi_n8__branch_10__data__0__anchor__in,
	input branch_15__Buffer_51__valid__0__anchor__in,
	input fork_17__branch_12__data__0__anchor__in,
	input fork_2__branch_7__ready__0__anchor__in,
	input [31 : 0] load_6__MC_A__data__0__anchor__in,
	input fork_16__branch_7__data__0__anchor__in,
	input [31 : 0] fork_4__branch_20__data__0__anchor__in,
	input icmp_0__fork_22__valid__0__anchor__in,
	input branch_19__sink_11__valid__0__anchor__in,
	input branch_17__sink_9__ready__0__anchor__in,
	input Buffer_54__phi_n7__ready__0__anchor__in,
	input branch_18__Buffer_53__ready__0__anchor__in,
	input [31 : 0] cst_3__add_11__data__0__anchor__in,
	input fork_16__branchC_24__data__0__anchor__in,
	input forkC_23__cst_1__ready__0__anchor__in,
	input forkC_28__branchC_27__data__0__anchor__in,
	input fork_14__branchC_22__ready__0__anchor__in,
	input [31 : 0] branch_3__phi_n6__data__0__anchor__in,
	input phi_n7__branch_9__ready__0__anchor__in,
	input MC_A__end_0__valid__0__anchor__in,
	input phi_n5__fork_4__ready__0__anchor__in,
	input branch_10__phi_n16__valid__0__anchor__in,
	input fork_10__branch_12__valid__0__anchor__in,
	input branchC_24__phiC_20__data__0__anchor__in,
	input forkC_23__branchC_22__valid__0__anchor__in,
	input fork_15__branch_4__ready__0__anchor__in,
	input MC_A__load_20__valid__0__anchor__in,
	input brCst_block3__fork_15__valid__0__anchor__in,
	input fork_18__branch_17__data__0__anchor__in,
	input brCst_block2__fork_14__data__0__anchor__in,
	input fork_16__branch_9__ready__0__anchor__in,
	input phiC_21__forkC_27__valid__0__anchor__in,
	input phi_8__fork_2__ready__0__anchor__in,
	input cst_2__icmp_9__ready__0__anchor__in,
	input add_17__load_20__ready__0__anchor__in,
	input fork_14__branch_1__data__0__anchor__in,
	input fork_18__branch_15__valid__0__anchor__in,
	input Buffer_58__fork_17__ready__0__anchor__in,
	input Buffer_53__phi_n8__ready__0__anchor__in,
	input phiC_22__forkC_28__data__0__anchor__in,
	input [31 : 0] phi_n3__store_1__data__0__anchor__in,
	input cst_7__MC_A__ready__0__anchor__in,
	input [30 : 0] branch_5__sink_5__data__0__anchor__in,
	input [31 : 0] fork_8__add_23__data__0__anchor__in,
	input fork_0__branch_0__valid__0__anchor__in,
	input branch_18__Buffer_53__valid__0__anchor__in,
	input fork_15__branch_6__data__0__anchor__in,
	input fork_19__branchC_27__data__0__anchor__in,
	input phi_n7__branch_9__valid__0__anchor__in,
	input [31 : 0] branch_14__phi_n12__data__0__anchor__in,
	input phiC_19__phi_8__data__0__anchor__in,
	input [30 : 0] fork_1__branch_6__data__0__anchor__in,
	input fork_8__add_17__valid__0__anchor__in,
	input [31 : 0] add_11__load_14__data__0__anchor__in,
	input fork_22__branch_0__valid__0__anchor__in,
	input fork_16__branch_7__ready__0__anchor__in,
	input phiC_18__phi_3__ready__0__anchor__in,
	input [31 : 0] cst_0__icmp_0__data__0__anchor__in,
	input branch_5__sink_5__valid__0__anchor__in,
	input phiC_21__forkC_27__data__0__anchor__in,
	input fork_16__branch_8__data__0__anchor__in,
	input Buffer_50__phi_n1__ready__0__anchor__in,
	input cst_8__MC_A__ready__0__anchor__in,
	input branchC_21__phiC_17__data__0__anchor__in,
	input branchC_25__phiC_21__data__0__anchor__in,
	input load_14__icmp_15__valid__0__anchor__in,
	input phi_n10__branch_16__valid__0__anchor__in,
	input fork_14__branch_2__ready__0__anchor__in,
	input branch_3__sink_3__valid__0__anchor__in,
	input phiC_19__phi_8__ready__0__anchor__in,
	input [31 : 0] cst_5__add_23__data__0__anchor__in,
	input load_14__icmp_15__ready__0__anchor__in,
	input fork_3__branch_19__valid__0__anchor__in,
	input [30 : 0] branch_19__Buffer_52__data__0__anchor__in,
	input branchC_24__phiC_22__valid__0__anchor__in,
	input [31 : 0] source_4__cst_5__data__0__anchor__in,
	input [31 : 0] fork_10__icmp_15__data__0__anchor__in,
	input forkC_27__branchC_26__data__0__anchor__in,
	input fork_17__branch_13__valid__0__anchor__in,
	input forkC_28__branchC_27__ready__0__anchor__in,
	input forkC_27__brCst_block6__ready__0__anchor__in,
	input [31 : 0] branch_16__sink_8__data__0__anchor__in,
	input Buffer_51__phi_8__valid__0__anchor__in,
	input [30 : 0] phi_n4__add_27__data__0__anchor__in,
	input forkC_23__cst_1__data__0__anchor__in,
	input icmp_9__fork_16__ready__0__anchor__in,
	input fork_15__branchC_23__ready__0__anchor__in,
	input fork_18__branch_18__ready__0__anchor__in,
	input fork_17__branchC_25__valid__0__anchor__in,
	input fork_10__icmp_15__ready__0__anchor__in,
	input [31 : 0] phi_n16__branch_14__data__0__anchor__in,
	input fork_19__branch_20__data__0__anchor__in,
	input forkC_27__brCst_block6__valid__0__anchor__in,
	input [31 : 0] branch_8__phi_n2__data__0__anchor__in,
	input fork_4__icmp_28__valid__0__anchor__in,
	input fork_16__branch_10__data__0__anchor__in,
	input branch_11__phi_n9__valid__0__anchor__in,
	input phiC_17__forkC_23__valid__0__anchor__in,
	input phi_n0__branch_2__valid__0__anchor__in,
	input MC_A__load_6__ready__0__anchor__in,
	input phi_n16__branch_14__valid__0__anchor__in,
	input branch_15__sink_7__ready__0__anchor__in,
	input [31 : 0] MC_A__load_20__data__0__anchor__in,
	input fork_4__branch_20__valid__0__anchor__in,
	input branch_1__sink_1__ready__0__anchor__in,
	input fork_14__branch_1__valid__0__anchor__in,
	input fork_15__branch_5__valid__0__anchor__in,
	input phi_n2__store_1__ready__0__anchor__in,
	input load_6__branch_3__ready__0__anchor__in,
	input icmp_28__fork_19__ready__0__anchor__in,
	input fork_14__branch_2__valid__0__anchor__in,
	input branchC_23__phiC_19__data__0__anchor__in,
	input cst_4__add_17__valid__0__anchor__in,
	input icmp_0__fork_22__ready__0__anchor__in,
	input add_27__fork_3__ready__0__anchor__in,
	input phi_n6__branch_8__valid__0__anchor__in,
	input [31 : 0] branch_12__phi_n10__data__0__anchor__in,
	input fork_16__branch_9__data__0__anchor__in,
	input brCst_block6__fork_18__data__0__anchor__in,
	input source_1__cst_2__data__0__anchor__in,
	input start_valid,
	input [31 : 0] branch_10__phi_n16__data__0__anchor__in,
	input fork_19__branchC_27__ready__0__anchor__in,
	input fork_22__branchC_21__data__0__anchor__in,
	input load_6__MC_A__valid__0__anchor__in,
	input n__fork_0__valid__0__anchor__in,
	input fork_17__branch_14__data__0__anchor__in,
	input [31 : 0] fork_3__icmp_28__data__0__anchor__in,
	input store_1__MC_A__valid__0__anchor__in,
	input [31 : 0] phi_n6__branch_8__data__0__anchor__in,
	input branchC_22__phiC_18__ready__0__anchor__in,
	input fork_15__branch_3__data__0__anchor__in,
	input [30 : 0] branch_17__sink_9__data__0__anchor__in,
	input [31 : 0] branch_8__phi_n14__data__0__anchor__in,
	input MC_A__load_14__ready__0__anchor__in,
	input Buffer_57__phiC_19__valid__0__anchor__in,
	input fork_17__branch_14__valid__0__anchor__in,
	input [31 : 0] phi_n12__branch_18__data__0__anchor__in,
	input phiC_19__phi_8__valid__0__anchor__in,
	input branch_1__phi_3__valid__0__anchor__in,
	input [30 : 0] branch_13__phi_n11__data__0__anchor__in,
	input branchC_23__phiC_19__valid__0__anchor__in,
	input branch_20__Buffer_50__ready__0__anchor__in,
	input [31 : 0] phi_n5__fork_4__data__0__anchor__in,
	input fork_17__branch_11__valid__0__anchor__in,
	input [31 : 0] phi_n0__branch_2__data__0__anchor__in,
	input Buffer_50__phi_n1__valid__0__anchor__in,
	input cst_2__icmp_9__valid__0__anchor__in,
	input cst_3__add_11__ready__0__anchor__in,
	input phi_n11__branch_17__ready__0__anchor__in,
	input [31 : 0] branch_6__phi_8__data__0__anchor__in,
	input fork_8__add_17__ready__0__anchor__in,
	input branch_10__phi_n16__ready__0__anchor__in,
	input [31 : 0] branch_20__sink_12__data__0__anchor__in,
	input Buffer_55__phi_n6__ready__0__anchor__in,
	input [31 : 0] load_14__icmp_15__data__0__anchor__in,
	input [31 : 0] branch_15__sink_7__data__0__anchor__in,
	input load_20__MC_A__valid__0__anchor__in,
	input [31 : 0] store_1__MC_A__data__0__anchor__in,
	input store_1__MC_A__valid__1__anchor__in,
	input branch_16__sink_8__valid__0__anchor__in,
	input [31 : 0] A_din1,
	input MC_A__load_14__valid__0__anchor__in,
	input branchC_25__phiC_22__valid__0__anchor__in,
	input phiC_23__ret_0__ready__0__anchor__in,
	input branchC_26__sink_15__valid__0__anchor__in,
	input branch_8__phi_n14__valid__0__anchor__in,
	input [30 : 0] fork_1__load_6__data__0__anchor__in,
	input load_14__MC_A__valid__0__anchor__in,
	input ret_0__end_0__data__0__anchor__in,
	input [30 : 0] fork_1__branch_5__data__0__anchor__in,
	input [30 : 0] branch_6__sink_6__data__0__anchor__in,
	input fork_17__branchC_25__data__0__anchor__in,
	input fork_8__add_23__ready__0__anchor__in,
	input fork_4__branch_20__ready__0__anchor__in,
	input phi_n15__branch_13__ready__0__anchor__in,
	input fork_15__branch_5__ready__0__anchor__in,
	input fork_1__branch_5__ready__0__anchor__in,
	input [30 : 0] branch_13__phi_n4__data__0__anchor__in,
	input branch_13__phi_n11__valid__0__anchor__in,
	input fork_18__branch_18__valid__0__anchor__in,
	input fork_17__branch_12__ready__0__anchor__in,
	input branchC_27__Buffer_56__valid__0__anchor__in,
	input [31 : 0] branch_7__phi_n3__data__0__anchor__in,
	input [31 : 0] branch_7__phi_n13__data__0__anchor__in,
	input icmp_9__fork_16__valid__0__anchor__in,
	input [31 : 0] fork_2__branch_7__data__0__anchor__in,
	input branch_16__Buffer_55__valid__0__anchor__in,
	input phi_n4__add_27__ready__0__anchor__in,
	input [31 : 0] branch_11__phi_n3__data__0__anchor__in,
	input branch_4__sink_4__valid__0__anchor__in,
	input branchC_23__sink_14__valid__0__anchor__in,
	input fork_9__branch_11__ready__0__anchor__in,
	input Buffer_57__phiC_19__ready__0__anchor__in,
	input forkC_23__brCst_block2__valid__0__anchor__in,
	input fork_19__branch_19__ready__0__anchor__in,
	input [31 : 0] source_3__cst_4__data__0__anchor__in,
	input [31 : 0] branch_14__phi_n5__data__0__anchor__in,
	input fork_15__branch_6__ready__0__anchor__in,
	input forkC_24__brCst_block3__ready__0__anchor__in,
	input phiC_19__branchC_24__data__0__anchor__in,
	input branch_13__phi_n11__ready__0__anchor__in,
	input cst_7__MC_A__valid__0__anchor__in,
	input [30 : 0] phi_3__fork_1__data__0__anchor__in,
	input phi_3__fork_1__valid__0__anchor__in,
	input fork_18__branch_17__ready__0__anchor__in,
	input cst_8__MC_A__valid__0__anchor__in,
	input branchC_27__phiC_23__ready__0__anchor__in,
	input branchC_26__sink_15__data__0__anchor__in,
	input fork_16__branch_10__valid__0__anchor__in,
	input [31 : 0] n_din,
	input branch_14__phi_n5__ready__0__anchor__in,
	input [31 : 0] fork_9__branch_11__data__0__anchor__in,
	input phi_n12__branch_18__valid__0__anchor__in,
	input branch_4__phi_n8__valid__0__anchor__in,
	input fork_16__branch_7__valid__0__anchor__in,
	input branchC_22__phiC_18__data__0__anchor__in,
	input branch_5__sink_5__ready__0__anchor__in,
	input [31 : 0] cst_7__MC_A__data__0__anchor__in,
	input source_1__cst_2__valid__0__anchor__in,
	input branch_9__phi_n15__valid__0__anchor__in,
	input cst_1__branch_1__data__0__anchor__in,
	input brCst_block3__fork_15__data__0__anchor__in,
	input branch_12__phi_n2__ready__0__anchor__in,
	input branch_11__phi_n9__ready__0__anchor__in,
	input branch_20__sink_12__ready__0__anchor__in,
	input phi_n9__fork_8__valid__0__anchor__in,
	input fork_19__branch_20__valid__0__anchor__in,
	input fork_18__branch_16__ready__0__anchor__in,
	input branch_6__phi_8__ready__0__anchor__in,
	input fork_3__icmp_28__ready__0__anchor__in,
	input branch_18__sink_10__valid__0__anchor__in,
	input fork_0__icmp_0__ready__0__anchor__in,
	input branchC_21__phiC_23__data__0__anchor__in,
	input fork_19__branch_20__ready__0__anchor__in,
	input [30 : 0] branch_17__Buffer_54__data__0__anchor__in,
	input phiC_18__forkC_24__valid__0__anchor__in,
	input branch_4__sink_4__ready__0__anchor__in,
	input [31 : 0] branch_2__phi_n1__data__0__anchor__in,
	input phi_n12__branch_18__ready__0__anchor__in,
	input branch_6__phi_8__valid__0__anchor__in,
	input branch_19__Buffer_52__valid__0__anchor__in,
	input forkC_27__brCst_block6__data__0__anchor__in,
	input branch_7__phi_n13__valid__0__anchor__in,
	input fork_2__branch_7__valid__0__anchor__in,
	input branchC_24__phiC_22__ready__0__anchor__in,
	input branchC_25__phiC_22__ready__0__anchor__in,
	input source_2__cst_3__ready__0__anchor__in,
	input Buffer_56__phiC_18__ready__0__anchor__in,
	input branch_8__phi_n14__ready__0__anchor__in,
	input start_0__branchC_21__ready__0__anchor__in,
	input add_17__load_20__valid__0__anchor__in,
	input [30 : 0] Buffer_54__phi_n7__data__0__anchor__in,
	input brCst_block3__fork_15__ready__0__anchor__in,
	input store_0__MC_A__ready__1__anchor__in,
	input Buffer_51__phi_8__ready__0__anchor__in,
	input load_6__MC_A__ready__0__anchor__in,
	input fork_18__branch_17__valid__0__anchor__in,
	input end_ready,
	input store_0__MC_A__valid__1__anchor__in,
	input cst_1__branch_1__valid__0__anchor__in,
	input branch_7__phi_n13__ready__0__anchor__in,
	input branchC_21__phiC_17__ready__0__anchor__in,
	input source_4__cst_5__valid__0__anchor__in,
	input [31 : 0] phi_n9__fork_8__data__0__anchor__in,
	input fork_16__branch_10__ready__0__anchor__in,
	input branch_15__sink_7__valid__0__anchor__in,
	input load_20__store_0__valid__0__anchor__in,
	input add_23__branch_15__ready__0__anchor__in,
	input store_0__MC_A__ready__0__anchor__in,
	input fork_14__branch_1__ready__0__anchor__in,
	input fork_17__branch_11__data__0__anchor__in,
	input branchC_26__Buffer_57__data__0__anchor__in,
	input fork_1__load_6__ready__0__anchor__in,
	input fork_18__branchC_26__valid__0__anchor__in,
	input forkC_28__cst_8__data__0__anchor__in,
	input branch_19__sink_11__ready__0__anchor__in,
	input [30 : 0] cst_6__add_27__data__0__anchor__in,
	input fork_9__add_11__valid__0__anchor__in,
	input branch_12__phi_n10__ready__0__anchor__in,
	input fork_15__branch_4__data__0__anchor__in,
	input fork_15__branch_3__ready__0__anchor__in,
	input brCst_block2__fork_14__ready__0__anchor__in,
	input [31 : 0] cst_8__MC_A__data__0__anchor__in,
	input branch_2__phi_n1__valid__0__anchor__in,
	input rst,
	input MC_A__end_0__ready__0__anchor__in,
	input branch_13__phi_n4__ready__0__anchor__in,
	input phi_n13__fork_9__valid__0__anchor__in,
	input branchC_24__phiC_22__data__0__anchor__in,
	input cst_4__add_17__ready__0__anchor__in,
	input Buffer_55__phi_n6__valid__0__anchor__in,
	input add_11__load_14__ready__0__anchor__in,
	input fork_8__store_0__ready__0__anchor__in,
	input start_in,
	input [31 : 0] branch_12__phi_n2__data__0__anchor__in,
	input [31 : 0] branch_0__phi_n0__data__0__anchor__in,
	input [31 : 0] fork_0__branch_0__data__0__anchor__in,
	input branch_17__Buffer_54__ready__0__anchor__in,
	input [31 : 0] phi_8__fork_2__data__0__anchor__in,
	input [31 : 0] source_2__cst_3__data__0__anchor__in,
	input [31 : 0] fork_10__branch_12__data__0__anchor__in,
	input forkC_28__branchC_27__valid__0__anchor__in,
	input fork_17__branchC_25__ready__0__anchor__in,
	input [31 : 0] MC_A__load_14__data__0__anchor__in,
	input cst_0__icmp_0__ready__0__anchor__in,
	input phiC_23__ret_0__data__0__anchor__in,
	input Buffer_52__phi_3__ready__0__anchor__in,
	input fork_15__branchC_23__data__0__anchor__in,
	input branchC_23__sink_14__ready__0__anchor__in,
	input branchC_25__phiC_22__data__0__anchor__in,
	input phi_n11__branch_17__valid__0__anchor__in,
	input fork_9__branch_11__valid__0__anchor__in,
	input fork_22__branchC_21__ready__0__anchor__in,
	input fork_1__branch_6__valid__0__anchor__in,
	input [30 : 0] fork_3__branch_19__data__0__anchor__in,
	input brCst_block6__fork_18__ready__0__anchor__in,
	input phi_n6__branch_8__ready__0__anchor__in,
	input [30 : 0] phi_n11__branch_17__data__0__anchor__in,
	input phi_n3__store_1__valid__0__anchor__in,
	input fork_14__branchC_22__data__0__anchor__in,
	input forkC_27__cst_7__valid__0__anchor__in,
	input branch_8__phi_n2__ready__0__anchor__in,
	input source_0__cst_0__ready__0__anchor__in,
	input branchC_27__Buffer_56__ready__0__anchor__in,
	input branch_10__phi_n5__valid__0__anchor__in,
	input icmp_15__Buffer_58__ready__0__anchor__in,
	input fork_9__add_11__ready__0__anchor__in,
	input branch_0__phi_n0__valid__0__anchor__in,
	input fork_18__branch_16__data__0__anchor__in,
	input branch_9__phi_n4__ready__0__anchor__in,
	input phiC_17__forkC_23__ready__0__anchor__in,
	input clk,
	input fork_2__icmp_9__ready__0__anchor__in,
	input source_1__cst_2__ready__0__anchor__in,
	input [30 : 0] branch_19__sink_11__data__0__anchor__in,
	input branch_16__Buffer_55__ready__0__anchor__in,
	input phiC_18__forkC_24__data__0__anchor__in,
	input source_5__cst_6__ready__0__anchor__in,
	input branchC_26__Buffer_57__ready__0__anchor__in,
	input branch_5__phi_n7__ready__0__anchor__in,
	input phiC_19__branchC_24__ready__0__anchor__in,
	input forkC_27__cst_7__data__0__anchor__in,
	input fork_10__icmp_15__valid__0__anchor__in,
	input branch_2__sink_2__valid__0__anchor__in,
	input branch_2__sink_2__ready__0__anchor__in,
	input phiC_22__forkC_28__ready__0__anchor__in,
	input forkC_28__cst_8__valid__0__anchor__in,
	input Buffer_56__phiC_18__valid__0__anchor__in,
	input [31 : 0] n__fork_0__data__0__anchor__in,
	input load_14__MC_A__ready__0__anchor__in,
	input [31 : 0] cst_2__icmp_9__data__0__anchor__in,
	input load_6__branch_3__valid__0__anchor__in,
	input fork_18__branch_18__data__0__anchor__in,
	input phiC_23__ret_0__valid__0__anchor__in,
	input fork_19__branch_19__valid__0__anchor__in,
	input [31 : 0] phi_n10__branch_16__data__0__anchor__in,
	input branch_12__phi_n10__valid__0__anchor__in,
	input fork_2__icmp_9__valid__0__anchor__in,
	input forkC_24__brCst_block3__valid__0__anchor__in,
	input branch_6__sink_6__ready__0__anchor__in,
	input Buffer_58__fork_17__valid__0__anchor__in,
	input [31 : 0] phi_n13__fork_9__data__0__anchor__in,
	input [31 : 0] Buffer_58__fork_17__data__0__anchor__in,
	input fork_16__branch_8__valid__0__anchor__in,
	input fork_15__branch_3__valid__0__anchor__in,
	input phiC_19__branchC_24__valid__0__anchor__in,
	input [31 : 0] fork_0__icmp_0__data__0__anchor__in,
	input phiC_18__phi_3__data__0__anchor__in,
	input [31 : 0] cst_4__add_17__data__0__anchor__in,
	input store_1__MC_A__ready__1__anchor__in,
	input branch_7__phi_n3__ready__0__anchor__in,
	input branch_9__phi_n15__ready__0__anchor__in,
	input [30 : 0] Buffer_52__phi_3__data__0__anchor__in,
	input phi_n15__branch_13__valid__0__anchor__in,
	input add_11__load_14__valid__0__anchor__in,
	input [31 : 0] load_14__MC_A__data__0__anchor__in,
	input Buffer_53__phi_n8__valid__0__anchor__in,
	input forkC_23__branchC_22__data__0__anchor__in,
	input start_0__branchC_21__valid__0__anchor__in,
	input [31 : 0] Buffer_50__phi_n1__data__0__anchor__in,
	input phi_n16__branch_14__ready__0__anchor__in,
	input [31 : 0] phi_n14__fork_10__data__0__anchor__in,
	input fork_17__branch_14__ready__0__anchor__in,
	input branchC_24__phiC_20__ready__0__anchor__in,
	input fork_17__branch_12__valid__0__anchor__in,
	input branch_1__sink_1__data__0__anchor__in,
	input branchC_23__phiC_19__ready__0__anchor__in,
	input phi_n1__branch_4__valid__0__anchor__in,
	input branch_0__sink_0__ready__0__anchor__in,
	input Buffer_56__phiC_18__data__0__anchor__in,
	input branchC_27__phiC_23__data__0__anchor__in,
	input [31 : 0] load_20__MC_A__data__0__anchor__in,
	input phiC_20__branchC_25__ready__0__anchor__in,
	input icmp_28__fork_19__data__0__anchor__in,
	input fork_15__branch_4__valid__0__anchor__in,
	input phi_n5__fork_4__valid__0__anchor__in,
	input [31 : 0] branch_18__sink_10__data__0__anchor__in,
	input [30 : 0] branch_9__phi_n15__data__0__anchor__in,
	input forkC_27__cst_7__ready__0__anchor__in,
	input fork_10__branch_12__ready__0__anchor__in,
	input store_0__MC_A__valid__0__anchor__in,
	input store_1__MC_A__ready__0__anchor__in,
	input branch_0__sink_0__valid__0__anchor__in,
	input source_3__cst_4__valid__0__anchor__in,
	input [31 : 0] branch_10__phi_n5__data__0__anchor__in,
	input phi_n2__store_1__valid__0__anchor__in,
	input fork_1__branch_5__valid__0__anchor__in,
	input [31 : 0] MC_A__load_6__data__0__anchor__in,
	input branch_17__Buffer_54__valid__0__anchor__in,
	input [31 : 0] store_0__MC_A__data__1__anchor__in,
	input Buffer_57__phiC_19__data__0__anchor__in,
	input [30 : 0] branch_9__phi_n4__data__0__anchor__in,
	input [31 : 0] branch_2__sink_2__data__0__anchor__in,
	input phi_n14__fork_10__ready__0__anchor__in,
	input fork_8__add_23__valid__0__anchor__in,
	input branchC_22__phiC_18__valid__0__anchor__in,
	input [31 : 0] load_20__store_0__data__0__anchor__in,
	input [31 : 0] fork_9__add_11__data__0__anchor__in,
	input branchC_21__phiC_23__valid__0__anchor__in,
	input fork_14__branchC_22__valid__0__anchor__in,
	input phi_n3__store_1__ready__0__anchor__in,
	input branch_4__phi_n8__ready__0__anchor__in,
	input branchC_25__phiC_21__ready__0__anchor__in,
	input phi_n1__branch_4__ready__0__anchor__in,
	input [30 : 0] phi_n15__branch_13__data__0__anchor__in,
	input forkC_27__branchC_26__valid__0__anchor__in,
	input fork_8__store_0__valid__0__anchor__in,
	input cst_6__add_27__ready__0__anchor__in,
	input phiC_18__forkC_24__ready__0__anchor__in,
	input branchC_27__phiC_23__valid__0__anchor__in,
	input fork_4__icmp_28__ready__0__anchor__in,
	input [31 : 0] add_17__load_20__data__0__anchor__in,
	input branchC_26__Buffer_57__valid__0__anchor__in,
	input cst_6__add_27__valid__0__anchor__in,
	input branch_10__phi_n5__ready__0__anchor__in,
	input Buffer_52__phi_3__valid__0__anchor__in,
	input branch_15__Buffer_51__ready__0__anchor__in,
	input [31 : 0] Buffer_51__phi_8__data__0__anchor__in,
	input cst_1__branch_1__ready__0__anchor__in,
	input Buffer_54__phi_n7__valid__0__anchor__in,
	input ret_0__end_0__ready__0__anchor__in,
	input cst_5__add_23__valid__0__anchor__in,
	input branch_7__phi_n3__valid__0__anchor__in,
	input branch_9__phi_n4__valid__0__anchor__in,
	input [31 : 0] branch_16__Buffer_55__data__0__anchor__in,
	input branchC_27__Buffer_56__data__0__anchor__in,
	input fork_14__branch_2__data__0__anchor__in,
	input phi_n0__branch_2__ready__0__anchor__in,
	input [31 : 0] store_1__MC_A__data__1__anchor__in,
	input [31 : 0] add_23__branch_15__data__0__anchor__in,
	input fork_16__branchC_24__ready__0__anchor__in,
	input [31 : 0] branch_11__phi_n9__data__0__anchor__in,
	input fork_1__branch_6__ready__0__anchor__in,
	input fork_17__branch_13__ready__0__anchor__in,
	input [31 : 0] A_din0,
	input [31 : 0] branch_0__sink_0__data__0__anchor__in,
	input branch_5__phi_n7__valid__0__anchor__in,
	input fork_22__branch_0__ready__0__anchor__in,
	input phi_n14__fork_10__valid__0__anchor__in,
	input source_2__cst_3__valid__0__anchor__in,
	input [31 : 0] load_6__branch_3__data__0__anchor__in,
	input [30 : 0] branch_1__phi_3__data__0__anchor__in,
	input icmp_9__fork_16__data__0__anchor__in,
	input branchC_24__phiC_20__valid__0__anchor__in,
	input phi_3__fork_1__ready__0__anchor__in,
	input branch_20__sink_12__valid__0__anchor__in,
	input [31 : 0] fork_2__icmp_9__data__0__anchor__in,
	input branchC_23__sink_14__data__0__anchor__in,
	input branch_19__Buffer_52__ready__0__anchor__in,
	input branch_14__phi_n12__valid__0__anchor__in,
	input fork_18__branch_15__data__0__anchor__in,
	input fork_0__icmp_0__valid__0__anchor__in,
	input forkC_24__brCst_block3__data__0__anchor__in,
	input cst_0__icmp_0__valid__0__anchor__in,
	input branchC_22__sink_13__ready__0__anchor__in,
	input branch_3__phi_n6__valid__0__anchor__in,
	input branch_20__Buffer_50__valid__0__anchor__in,
	input [31 : 0] branch_4__sink_4__data__0__anchor__in,
	input icmp_0__fork_22__data__0__anchor__in,
	input fork_15__branch_5__data__0__anchor__in,
	input branch_11__phi_n3__valid__0__anchor__in,
	input MC_A__end_0__data__0__anchor__in,
	input [1 : 0] source_0__cst_0__data__0__anchor__in,
	input add_23__branch_15__valid__0__anchor__in,
	input brCst_block2__fork_14__valid__0__anchor__in,
	input [31 : 0] phi_n1__branch_4__data__0__anchor__in,
	input branch_2__phi_n1__ready__0__anchor__in,
	input branch_14__phi_n12__ready__0__anchor__in,
	input branch_6__sink_6__valid__0__anchor__in,
	input brCst_block6__fork_18__valid__0__anchor__in,
	input add_27__fork_3__valid__0__anchor__in,
	input phiC_20__branchC_25__data__0__anchor__in,
	input branch_3__sink_3__ready__0__anchor__in,
	input icmp_28__fork_19__valid__0__anchor__in,
	input phiC_20__branchC_25__valid__0__anchor__in,
	input branchC_26__sink_15__ready__0__anchor__in,
	input source_5__cst_6__data__0__anchor__in,
	input n__fork_0__ready__0__anchor__in,
	input fork_15__branchC_23__valid__0__anchor__in,
	input [31 : 0] branch_18__Buffer_53__data__0__anchor__in,
	input fork_22__branchC_21__valid__0__anchor__in,
	input fork_3__branch_19__ready__0__anchor__in,
	input [31 : 0] fork_4__icmp_28__data__0__anchor__in,
	input fork_17__branch_13__data__0__anchor__in,
	input branchC_22__sink_13__data__0__anchor__in,
	input branch_0__phi_n0__ready__0__anchor__in,
	input load_20__store_0__ready__0__anchor__in,
	input phiC_17__forkC_23__data__0__anchor__in,
	input branchC_22__sink_13__valid__0__anchor__in,
	input fork_3__icmp_28__valid__0__anchor__in,
	input fork_18__branchC_26__ready__0__anchor__in,
	input start_0__branchC_21__data__0__anchor__in,
	input phiC_18__phi_3__valid__0__anchor__in,
	input [31 : 0] branch_4__phi_n8__data__0__anchor__in,
	input fork_0__branch_0__ready__0__anchor__in,
	input source_0__cst_0__valid__0__anchor__in,
	input branchC_21__phiC_17__valid__0__anchor__in,
	input fork_19__branch_19__data__0__anchor__in,
	input source_5__cst_6__valid__0__anchor__in,
	input icmp_15__Buffer_58__valid__0__anchor__in,
	input MC_A__load_6__valid__0__anchor__in,
	input branch_14__phi_n5__valid__0__anchor__in,
	input branch_16__sink_8__ready__0__anchor__in,
	input cst_3__add_11__valid__0__anchor__in,
	input branch_1__sink_1__valid__0__anchor__in,
	input [31 : 0] icmp_15__Buffer_58__data__0__anchor__in,
	input forkC_24__branchC_23__ready__0__anchor__in,
	input cst_5__add_23__ready__0__anchor__in,
	input [31 : 0] Buffer_53__phi_n8__data__0__anchor__in,
	input [31 : 0] branch_3__sink_3__data__0__anchor__in,
	input fork_16__branch_8__ready__0__anchor__in,
	input forkC_24__branchC_23__valid__0__anchor__in,
	input forkC_23__brCst_block2__data__0__anchor__in,
	input fork_18__branch_15__ready__0__anchor__in,
	input fork_17__branch_11__ready__0__anchor__in,
	input source_4__cst_5__ready__0__anchor__in,
	input fork_16__branch_9__valid__0__anchor__in,
	input fork_19__branchC_27__valid__0__anchor__in,
	input load_20__MC_A__ready__0__anchor__in,
	input [31 : 0] phi_n2__store_1__data__0__anchor__in,
	input branchC_25__phiC_21__valid__0__anchor__in,
	input phi_n13__fork_9__ready__0__anchor__in,
	input fork_22__branch_0__data__0__anchor__in,
	input phi_n8__branch_10__valid__0__anchor__in,
	input [31 : 0] branch_15__Buffer_51__data__0__anchor__in,
	input phi_n9__fork_8__ready__0__anchor__in,
	input [30 : 0] branch_5__phi_n7__data__0__anchor__in,
	input source_3__cst_4__ready__0__anchor__in,
	input branchC_21__phiC_23__ready__0__anchor__in,
	input branch_11__phi_n3__ready__0__anchor__in,
	input n_valid_in,
	input phiC_21__forkC_27__ready__0__anchor__in,
	input fork_1__load_6__valid__0__anchor__in,
	input branch_18__sink_10__ready__0__anchor__in,
	input branch_13__phi_n4__valid__0__anchor__in,
	input [30 : 0] phi_n7__branch_9__data__0__anchor__in,
	input MC_A__load_20__ready__0__anchor__in,
	input [31 : 0] branch_20__Buffer_50__data__0__anchor__in,
	input phi_n4__add_27__valid__0__anchor__in,
	input forkC_24__branchC_23__data__0__anchor__in,
	input fork_16__branchC_24__valid__0__anchor__in,
	input ret_0__end_0__valid__0__anchor__in,
	input forkC_23__cst_1__valid__0__anchor__in,
	input [30 : 0] add_27__fork_3__data__0__anchor__in,
	input [31 : 0] store_0__MC_A__data__0__anchor__in,
	input branch_12__phi_n2__valid__0__anchor__in,
	input phiC_22__forkC_28__valid__0__anchor__in,
	input phi_n8__branch_10__ready__0__anchor__in,
	input fork_18__branchC_26__data__0__anchor__in,
	input branch_17__sink_9__valid__0__anchor__in,
	input phi_8__fork_2__valid__0__anchor__in,
	output A_ce1,
	output fork_9__branch_11__valid__0__anchor__out,
	output phi_n7__branch_9__ready__0__anchor__out,
	output [30 : 0] phi_3__fork_1__data__0__anchor__out,
	output branchC_27__phiC_23__valid__0__anchor__out,
	output [31 : 0] branch_2__phi_n1__data__0__anchor__out,
	output phiC_21__forkC_27__ready__0__anchor__out,
	output [31 : 0] cst_8__MC_A__data__0__anchor__out,
	output [31 : 0] branch_3__sink_3__data__0__anchor__out,
	output [31 : 0] branch_18__sink_10__data__0__anchor__out,
	output load_6__branch_3__valid__0__anchor__out,
	output branchC_24__phiC_22__valid__0__anchor__out,
	output [31 : 0] branch_11__phi_n9__data__0__anchor__out,
	output Buffer_52__phi_3__valid__0__anchor__out,
	output phi_n10__branch_16__ready__0__anchor__out,
	output branch_1__sink_1__data__0__anchor__out,
	output fork_1__branch_5__ready__0__anchor__out,
	output fork_9__add_11__valid__0__anchor__out,
	output branchC_22__phiC_18__valid__0__anchor__out,
	output fork_3__icmp_28__valid__0__anchor__out,
	output branchC_26__sink_15__ready__0__anchor__out,
	output fork_16__branch_9__data__0__anchor__out,
	output branch_14__phi_n12__ready__0__anchor__out,
	output branch_20__sink_12__ready__0__anchor__out,
	output branch_18__sink_10__ready__0__anchor__out,
	output forkC_23__brCst_block2__ready__0__anchor__out,
	output phiC_18__phi_3__data__0__anchor__out,
	output source_5__cst_6__data__0__anchor__out,
	output fork_22__branchC_21__ready__0__anchor__out,
	output store_1__MC_A__valid__0__anchor__out,
	output fork_8__add_17__ready__0__anchor__out,
	output branch_14__phi_n5__valid__0__anchor__out,
	output brCst_block3__fork_15__ready__0__anchor__out,
	output store_1__MC_A__ready__1__anchor__out,
	output [31 : 0] branch_6__phi_8__data__0__anchor__out,
	output fork_17__branchC_25__data__0__anchor__out,
	output branchC_27__Buffer_56__ready__0__anchor__out,
	output [31 : 0] cst_5__add_23__data__0__anchor__out,
	output fork_16__branch_10__ready__0__anchor__out,
	output branchC_21__phiC_23__data__0__anchor__out,
	output branch_15__Buffer_51__ready__0__anchor__out,
	output branchC_25__phiC_21__data__0__anchor__out,
	output [31 : 0] load_6__branch_3__data__0__anchor__out,
	output fork_19__branch_19__data__0__anchor__out,
	output forkC_27__brCst_block6__ready__0__anchor__out,
	output phi_n6__branch_8__valid__0__anchor__out,
	output brCst_block3__fork_15__valid__0__anchor__out,
	output icmp_9__fork_16__data__0__anchor__out,
	output branch_12__phi_n2__ready__0__anchor__out,
	output branchC_23__sink_14__valid__0__anchor__out,
	output phiC_22__forkC_28__valid__0__anchor__out,
	output [31 : 0] Buffer_58__fork_17__data__0__anchor__out,
	output fork_18__branch_15__valid__0__anchor__out,
	output fork_14__branchC_22__data__0__anchor__out,
	output fork_3__branch_19__ready__0__anchor__out,
	output fork_17__branch_11__data__0__anchor__out,
	output branchC_25__phiC_22__ready__0__anchor__out,
	output [31 : 0] branch_10__phi_n16__data__0__anchor__out,
	output start_0__branchC_21__valid__0__anchor__out,
	output branch_13__phi_n4__valid__0__anchor__out,
	output [31 : 0] source_3__cst_4__data__0__anchor__out,
	output forkC_23__cst_1__valid__0__anchor__out,
	output branchC_21__phiC_23__ready__0__anchor__out,
	output branch_16__Buffer_55__ready__0__anchor__out,
	output add_17__load_20__ready__0__anchor__out,
	output fork_14__branch_2__valid__0__anchor__out,
	output Buffer_57__phiC_19__valid__0__anchor__out,
	output phi_n0__branch_2__valid__0__anchor__out,
	output branch_7__phi_n3__valid__0__anchor__out,
	output icmp_0__fork_22__valid__0__anchor__out,
	output fork_17__branchC_25__ready__0__anchor__out,
	output store_0__MC_A__ready__0__anchor__out,
	output phi_3__fork_1__ready__0__anchor__out,
	output branch_13__phi_n4__ready__0__anchor__out,
	output [31 : 0] branch_16__sink_8__data__0__anchor__out,
	output n__fork_0__valid__0__anchor__out,
	output start_0__branchC_21__data__0__anchor__out,
	output forkC_23__brCst_block2__valid__0__anchor__out,
	output add_11__load_14__ready__0__anchor__out,
	output fork_16__branchC_24__ready__0__anchor__out,
	output [31 : 0] phi_n0__branch_2__data__0__anchor__out,
	output fork_1__branch_5__valid__0__anchor__out,
	output branch_10__phi_n16__ready__0__anchor__out,
	output fork_1__load_6__ready__0__anchor__out,
	output fork_16__branch_7__valid__0__anchor__out,
	output [31 : 0] phi_n3__store_1__data__0__anchor__out,
	output phiC_19__phi_8__data__0__anchor__out,
	output Buffer_57__phiC_19__ready__0__anchor__out,
	output [31 : 0] phi_n14__fork_10__data__0__anchor__out,
	output fork_0__branch_0__ready__0__anchor__out,
	output phi_n1__branch_4__ready__0__anchor__out,
	output [31 : 0] load_14__MC_A__data__0__anchor__out,
	output phiC_19__branchC_24__valid__0__anchor__out,
	output phi_n2__store_1__ready__0__anchor__out,
	output [30 : 0] phi_n11__branch_17__data__0__anchor__out,
	output source_1__cst_2__data__0__anchor__out,
	output [31 : 0] branch_11__phi_n3__data__0__anchor__out,
	output fork_15__branch_3__ready__0__anchor__out,
	output MC_A__end_0__ready__0__anchor__out,
	output [31 : 0] branch_8__phi_n14__data__0__anchor__out,
	output [30 : 0] Buffer_54__phi_n7__data__0__anchor__out,
	output branch_17__Buffer_54__ready__0__anchor__out,
	output branch_12__phi_n10__valid__0__anchor__out,
	output [31 : 0] store_0__MC_A__data__1__anchor__out,
	output [31 : 0] branch_8__phi_n2__data__0__anchor__out,
	output [31 : 0] add_11__load_14__data__0__anchor__out,
	output [30 : 0] branch_13__phi_n11__data__0__anchor__out,
	output branch_16__sink_8__valid__0__anchor__out,
	output add_11__load_14__valid__0__anchor__out,
	output cst_6__add_27__valid__0__anchor__out,
	output fork_0__branch_0__valid__0__anchor__out,
	output fork_15__branch_6__data__0__anchor__out,
	output [30 : 0] branch_9__phi_n4__data__0__anchor__out,
	output Buffer_50__phi_n1__ready__0__anchor__out,
	output branchC_24__phiC_20__valid__0__anchor__out,
	output phiC_18__forkC_24__valid__0__anchor__out,
	output load_20__store_0__valid__0__anchor__out,
	output Buffer_55__phi_n6__valid__0__anchor__out,
	output Buffer_51__phi_8__ready__0__anchor__out,
	output branch_7__phi_n13__valid__0__anchor__out,
	output load_20__store_0__ready__0__anchor__out,
	output [30 : 0] branch_5__sink_5__data__0__anchor__out,
	output brCst_block6__fork_18__valid__0__anchor__out,
	output load_20__MC_A__valid__0__anchor__out,
	output source_3__cst_4__valid__0__anchor__out,
	output phi_n2__store_1__valid__0__anchor__out,
	output icmp_28__fork_19__valid__0__anchor__out,
	output source_5__cst_6__valid__0__anchor__out,
	output branch_5__sink_5__ready__0__anchor__out,
	output [31 : 0] Buffer_50__phi_n1__data__0__anchor__out,
	output fork_15__branch_5__data__0__anchor__out,
	output phi_n15__branch_13__valid__0__anchor__out,
	output fork_18__branch_15__ready__0__anchor__out,
	output [31 : 0] fork_2__icmp_9__data__0__anchor__out,
	output [31 : 0] A_address1,
	output phiC_18__phi_3__valid__0__anchor__out,
	output forkC_28__cst_8__data__0__anchor__out,
	output phiC_21__forkC_27__valid__0__anchor__out,
	output [31 : 0] phi_n6__branch_8__data__0__anchor__out,
	output branchC_25__phiC_22__data__0__anchor__out,
	output fork_18__branchC_26__data__0__anchor__out,
	output [31 : 0] fork_8__add_17__data__0__anchor__out,
	output MC_A__load_6__ready__0__anchor__out,
	output branch_0__phi_n0__ready__0__anchor__out,
	output phi_n0__branch_2__ready__0__anchor__out,
	output phiC_18__phi_3__ready__0__anchor__out,
	output fork_18__branch_17__data__0__anchor__out,
	output icmp_9__fork_16__ready__0__anchor__out,
	output [31 : 0] MC_A__load_6__data__0__anchor__out,
	output [31 : 0] MC_A__load_14__data__0__anchor__out,
	output source_0__cst_0__valid__0__anchor__out,
	output branch_14__phi_n5__ready__0__anchor__out,
	output phiC_23__ret_0__data__0__anchor__out,
	output cst_1__branch_1__data__0__anchor__out,
	output fork_14__branch_2__data__0__anchor__out,
	output [30 : 0] branch_1__phi_3__data__0__anchor__out,
	output Buffer_53__phi_n8__valid__0__anchor__out,
	output fork_16__branch_9__valid__0__anchor__out,
	output branch_0__phi_n0__valid__0__anchor__out,
	output fork_8__add_23__ready__0__anchor__out,
	output fork_10__icmp_15__ready__0__anchor__out,
	output phiC_19__branchC_24__ready__0__anchor__out,
	output branchC_23__phiC_19__data__0__anchor__out,
	output fork_4__icmp_28__ready__0__anchor__out,
	output phiC_19__phi_8__valid__0__anchor__out,
	output icmp_9__fork_16__valid__0__anchor__out,
	output fork_18__branch_18__data__0__anchor__out,
	output phi_8__fork_2__ready__0__anchor__out,
	output fork_18__branch_17__ready__0__anchor__out,
	output branch_8__phi_n2__ready__0__anchor__out,
	output fork_14__branch_2__ready__0__anchor__out,
	output [31 : 0] fork_4__icmp_28__data__0__anchor__out,
	output [31 : 0] phi_n12__branch_18__data__0__anchor__out,
	output branch_11__phi_n9__valid__0__anchor__out,
	output icmp_28__fork_19__data__0__anchor__out,
	output fork_17__branch_11__ready__0__anchor__out,
	output fork_19__branch_19__ready__0__anchor__out,
	output branchC_24__phiC_20__data__0__anchor__out,
	output fork_22__branchC_21__data__0__anchor__out,
	output phi_n8__branch_10__valid__0__anchor__out,
	output load_14__icmp_15__valid__0__anchor__out,
	output branch_9__phi_n4__valid__0__anchor__out,
	output forkC_27__cst_7__ready__0__anchor__out,
	output fork_8__add_23__valid__0__anchor__out,
	output fork_16__branchC_24__data__0__anchor__out,
	output Buffer_56__phiC_18__valid__0__anchor__out,
	output [31 : 0] fork_8__add_23__data__0__anchor__out,
	output forkC_27__branchC_26__ready__0__anchor__out,
	output branchC_26__Buffer_57__ready__0__anchor__out,
	output fork_17__branch_13__ready__0__anchor__out,
	output [30 : 0] branch_17__Buffer_54__data__0__anchor__out,
	output end_out,
	output branch_6__sink_6__ready__0__anchor__out,
	output branchC_27__phiC_23__ready__0__anchor__out,
	output [30 : 0] branch_19__sink_11__data__0__anchor__out,
	output fork_19__branch_19__valid__0__anchor__out,
	output [31 : 0] branch_3__phi_n6__data__0__anchor__out,
	output [31 : 0] branch_7__phi_n3__data__0__anchor__out,
	output branch_19__Buffer_52__valid__0__anchor__out,
	output source_0__cst_0__ready__0__anchor__out,
	output branchC_22__phiC_18__data__0__anchor__out,
	output phi_3__fork_1__valid__0__anchor__out,
	output forkC_24__branchC_23__ready__0__anchor__out,
	output load_6__MC_A__valid__0__anchor__out,
	output branch_12__phi_n2__valid__0__anchor__out,
	output load_20__MC_A__ready__0__anchor__out,
	output [31 : 0] phi_n5__fork_4__data__0__anchor__out,
	output branch_5__phi_n7__ready__0__anchor__out,
	output [31 : 0] branch_12__phi_n10__data__0__anchor__out,
	output fork_17__branch_14__valid__0__anchor__out,
	output fork_14__branch_1__ready__0__anchor__out,
	output cst_6__add_27__ready__0__anchor__out,
	output branch_0__sink_0__ready__0__anchor__out,
	output branch_19__sink_11__ready__0__anchor__out,
	output [31 : 0] fork_10__branch_12__data__0__anchor__out,
	output branch_0__sink_0__valid__0__anchor__out,
	output fork_15__branchC_23__ready__0__anchor__out,
	output Buffer_51__phi_8__valid__0__anchor__out,
	output [31 : 0] fork_0__icmp_0__data__0__anchor__out,
	output fork_16__branch_8__data__0__anchor__out,
	output [31 : 0] source_2__cst_3__data__0__anchor__out,
	output [31 : 0] add_17__load_20__data__0__anchor__out,
	output source_3__cst_4__ready__0__anchor__out,
	output branchC_23__sink_14__ready__0__anchor__out,
	output icmp_0__fork_22__ready__0__anchor__out,
	output forkC_27__branchC_26__valid__0__anchor__out,
	output source_4__cst_5__valid__0__anchor__out,
	output ret_0__end_0__valid__0__anchor__out,
	output phi_n13__fork_9__ready__0__anchor__out,
	output branch_9__phi_n15__ready__0__anchor__out,
	output branch_2__phi_n1__valid__0__anchor__out,
	output cst_3__add_11__valid__0__anchor__out,
	output source_5__cst_6__ready__0__anchor__out,
	output Buffer_56__phiC_18__data__0__anchor__out,
	output phi_n13__fork_9__valid__0__anchor__out,
	output branchC_22__phiC_18__ready__0__anchor__out,
	output branch_11__phi_n9__ready__0__anchor__out,
	output branch_4__sink_4__ready__0__anchor__out,
	output [31 : 0] branch_12__phi_n2__data__0__anchor__out,
	output fork_18__branch_16__ready__0__anchor__out,
	output phi_n10__branch_16__valid__0__anchor__out,
	output branch_4__phi_n8__ready__0__anchor__out,
	output phi_n4__add_27__valid__0__anchor__out,
	output branch_11__phi_n3__ready__0__anchor__out,
	output branchC_21__phiC_23__valid__0__anchor__out,
	output branch_7__phi_n13__ready__0__anchor__out,
	output cst_7__MC_A__ready__0__anchor__out,
	output fork_17__branchC_25__valid__0__anchor__out,
	output fork_19__branchC_27__valid__0__anchor__out,
	output fork_8__add_17__valid__0__anchor__out,
	output [31 : 0] fork_9__add_11__data__0__anchor__out,
	output [31 : 0] load_14__icmp_15__data__0__anchor__out,
	output fork_16__branch_7__ready__0__anchor__out,
	output fork_18__branch_15__data__0__anchor__out,
	output [31 : 0] branch_15__Buffer_51__data__0__anchor__out,
	output branchC_21__phiC_17__valid__0__anchor__out,
	output add_17__load_20__valid__0__anchor__out,
	output phi_n1__branch_4__valid__0__anchor__out,
	output fork_19__branch_20__ready__0__anchor__out,
	output [31 : 0] branch_20__sink_12__data__0__anchor__out,
	output load_6__MC_A__ready__0__anchor__out,
	output branch_13__phi_n11__ready__0__anchor__out,
	output fork_2__branch_7__valid__0__anchor__out,
	output branch_15__Buffer_51__valid__0__anchor__out,
	output [30 : 0] branch_5__phi_n7__data__0__anchor__out,
	output phiC_23__ret_0__valid__0__anchor__out,
	output [31 : 0] branch_2__sink_2__data__0__anchor__out,
	output fork_18__branch_17__valid__0__anchor__out,
	output fork_1__branch_6__ready__0__anchor__out,
	output cst_4__add_17__valid__0__anchor__out,
	output branch_9__phi_n4__ready__0__anchor__out,
	output branch_18__Buffer_53__valid__0__anchor__out,
	output fork_19__branchC_27__data__0__anchor__out,
	output forkC_23__branchC_22__valid__0__anchor__out,
	output [31 : 0] Buffer_55__phi_n6__data__0__anchor__out,
	output branchC_26__sink_15__valid__0__anchor__out,
	output fork_2__icmp_9__ready__0__anchor__out,
	output fork_4__icmp_28__valid__0__anchor__out,
	output branchC_27__phiC_23__data__0__anchor__out,
	output brCst_block3__fork_15__data__0__anchor__out,
	output branch_10__phi_n5__ready__0__anchor__out,
	output branchC_22__sink_13__data__0__anchor__out,
	output branchC_22__sink_13__valid__0__anchor__out,
	output forkC_28__branchC_27__ready__0__anchor__out,
	output fork_8__store_0__ready__0__anchor__out,
	output branch_17__sink_9__valid__0__anchor__out,
	output phiC_18__forkC_24__ready__0__anchor__out,
	output ret_0__end_0__ready__0__anchor__out,
	output load_6__branch_3__ready__0__anchor__out,
	output fork_16__branch_10__data__0__anchor__out,
	output fork_22__branchC_21__valid__0__anchor__out,
	output branch_13__phi_n11__valid__0__anchor__out,
	output phiC_20__branchC_25__ready__0__anchor__out,
	output fork_19__branch_20__valid__0__anchor__out,
	output [31 : 0] phi_8__fork_2__data__0__anchor__out,
	output brCst_block2__fork_14__ready__0__anchor__out,
	output branch_11__phi_n3__valid__0__anchor__out,
	output [31 : 0] cst_0__icmp_0__data__0__anchor__out,
	output cst_0__icmp_0__ready__0__anchor__out,
	output forkC_23__cst_1__ready__0__anchor__out,
	output fork_0__icmp_0__ready__0__anchor__out,
	output forkC_24__brCst_block3__valid__0__anchor__out,
	output branch_6__phi_8__valid__0__anchor__out,
	output [31 : 0] A_address0,
	output MC_A__end_0__valid__0__anchor__out,
	output phi_n16__branch_14__ready__0__anchor__out,
	output forkC_28__branchC_27__data__0__anchor__out,
	output fork_15__branch_4__data__0__anchor__out,
	output fork_17__branch_14__ready__0__anchor__out,
	output branchC_25__phiC_21__valid__0__anchor__out,
	output branchC_27__Buffer_56__valid__0__anchor__out,
	output Buffer_57__phiC_19__data__0__anchor__out,
	output phi_n6__branch_8__ready__0__anchor__out,
	output branch_3__phi_n6__ready__0__anchor__out,
	output fork_15__branch_4__valid__0__anchor__out,
	output branch_18__sink_10__valid__0__anchor__out,
	output branch_1__phi_3__ready__0__anchor__out,
	output branchC_27__Buffer_56__data__0__anchor__out,
	output [30 : 0] branch_13__phi_n4__data__0__anchor__out,
	output phiC_17__forkC_23__ready__0__anchor__out,
	output fork_16__branch_8__valid__0__anchor__out,
	output [30 : 0] branch_17__sink_9__data__0__anchor__out,
	output icmp_15__Buffer_58__ready__0__anchor__out,
	output store_0__MC_A__ready__1__anchor__out,
	output brCst_block2__fork_14__data__0__anchor__out,
	output [31 : 0] cst_3__add_11__data__0__anchor__out,
	output [31 : 0] fork_0__branch_0__data__0__anchor__out,
	output fork_15__branch_5__valid__0__anchor__out,
	output fork_15__branch_6__ready__0__anchor__out,
	output phi_n3__store_1__valid__0__anchor__out,
	output [30 : 0] branch_6__sink_6__data__0__anchor__out,
	output [30 : 0] fork_1__load_6__data__0__anchor__out,
	output branch_20__Buffer_50__valid__0__anchor__out,
	output fork_22__branch_0__data__0__anchor__out,
	output fork_17__branch_12__ready__0__anchor__out,
	output cst_2__icmp_9__valid__0__anchor__out,
	output cst_4__add_17__ready__0__anchor__out,
	output fork_10__icmp_15__valid__0__anchor__out,
	output phi_n5__fork_4__ready__0__anchor__out,
	output branch_1__phi_3__valid__0__anchor__out,
	output A_ce0,
	output branch_10__phi_n16__valid__0__anchor__out,
	output [1 : 0] source_0__cst_0__data__0__anchor__out,
	output fork_14__branch_1__data__0__anchor__out,
	output fork_4__branch_20__ready__0__anchor__out,
	output fork_15__branch_5__ready__0__anchor__out,
	output branch_10__phi_n5__valid__0__anchor__out,
	output phiC_20__branchC_25__data__0__anchor__out,
	output [31 : 0] branch_10__phi_n5__data__0__anchor__out,
	output [31 : 0] cst_7__MC_A__data__0__anchor__out,
	output branch_2__phi_n1__ready__0__anchor__out,
	output fork_22__branch_0__valid__0__anchor__out,
	output branchC_23__phiC_19__valid__0__anchor__out,
	output [31 : 0] add_23__branch_15__data__0__anchor__out,
	output fork_18__branchC_26__ready__0__anchor__out,
	output n__fork_0__ready__0__anchor__out,
	output Buffer_58__fork_17__ready__0__anchor__out,
	output branch_17__sink_9__ready__0__anchor__out,
	output [31 : 0] load_20__store_0__data__0__anchor__out,
	output fork_4__branch_20__valid__0__anchor__out,
	output branchC_26__Buffer_57__data__0__anchor__out,
	output forkC_28__cst_8__valid__0__anchor__out,
	output [31 : 0] phi_n1__branch_4__data__0__anchor__out,
	output [31 : 0] source_4__cst_5__data__0__anchor__out,
	output Buffer_52__phi_3__ready__0__anchor__out,
	output branch_15__sink_7__ready__0__anchor__out,
	output [30 : 0] phi_n7__branch_9__data__0__anchor__out,
	output forkC_23__branchC_22__ready__0__anchor__out,
	output fork_16__branch_7__data__0__anchor__out,
	output fork_15__branch_3__valid__0__anchor__out,
	output fork_19__branchC_27__ready__0__anchor__out,
	output A_we0,
	output phi_n9__fork_8__ready__0__anchor__out,
	output [31 : 0] branch_4__sink_4__data__0__anchor__out,
	output fork_15__branch_4__ready__0__anchor__out,
	output fork_14__branchC_22__valid__0__anchor__out,
	output fork_16__branch_9__ready__0__anchor__out,
	output fork_2__icmp_9__valid__0__anchor__out,
	output [31 : 0] fork_9__branch_11__data__0__anchor__out,
	output forkC_23__brCst_block2__data__0__anchor__out,
	output branchC_24__phiC_22__ready__0__anchor__out,
	output MC_A__load_14__valid__0__anchor__out,
	output branch_3__sink_3__ready__0__anchor__out,
	output [31 : 0] icmp_15__Buffer_58__data__0__anchor__out,
	output phi_n4__add_27__ready__0__anchor__out,
	output store_0__MC_A__valid__0__anchor__out,
	output branch_6__phi_8__ready__0__anchor__out,
	output [31 : 0] Buffer_51__phi_8__data__0__anchor__out,
	output cst_1__branch_1__valid__0__anchor__out,
	output load_14__icmp_15__ready__0__anchor__out,
	output ret_0__end_0__data__0__anchor__out,
	output fork_3__icmp_28__ready__0__anchor__out,
	output branch_14__phi_n12__valid__0__anchor__out,
	output [31 : 0] branch_20__Buffer_50__data__0__anchor__out,
	output Buffer_54__phi_n7__ready__0__anchor__out,
	output phiC_22__forkC_28__ready__0__anchor__out,
	output add_27__fork_3__valid__0__anchor__out,
	output phi_n3__store_1__ready__0__anchor__out,
	output forkC_28__cst_8__ready__0__anchor__out,
	output [31 : 0] phi_n8__branch_10__data__0__anchor__out,
	output branch_2__sink_2__valid__0__anchor__out,
	output source_4__cst_5__ready__0__anchor__out,
	output add_27__fork_3__ready__0__anchor__out,
	output Buffer_58__fork_17__valid__0__anchor__out,
	output branchC_21__phiC_17__data__0__anchor__out,
	output [31 : 0] fork_2__branch_7__data__0__anchor__out,
	output MC_A__load_14__ready__0__anchor__out,
	output forkC_24__brCst_block3__data__0__anchor__out,
	output branch_2__sink_2__ready__0__anchor__out,
	output branch_8__phi_n2__valid__0__anchor__out,
	output phiC_22__forkC_28__data__0__anchor__out,
	output start_ready,
	output Buffer_50__phi_n1__valid__0__anchor__out,
	output branch_12__phi_n10__ready__0__anchor__out,
	output MC_A__load_20__valid__0__anchor__out,
	output [31 : 0] cst_4__add_17__data__0__anchor__out,
	output [30 : 0] branch_19__Buffer_52__data__0__anchor__out,
	output phi_n12__branch_18__ready__0__anchor__out,
	output load_14__MC_A__valid__0__anchor__out,
	output forkC_27__brCst_block6__valid__0__anchor__out,
	output branchC_23__phiC_19__ready__0__anchor__out,
	output add_23__branch_15__valid__0__anchor__out,
	output cst_1__branch_1__ready__0__anchor__out,
	output branchC_26__Buffer_57__valid__0__anchor__out,
	output phi_8__fork_2__valid__0__anchor__out,
	output Buffer_55__phi_n6__ready__0__anchor__out,
	output source_2__cst_3__valid__0__anchor__out,
	output branch_1__sink_1__valid__0__anchor__out,
	output [31 : 0] branch_0__phi_n0__data__0__anchor__out,
	output [31 : 0] phi_n9__fork_8__data__0__anchor__out,
	output [31 : 0] branch_4__phi_n8__data__0__anchor__out,
	output fork_16__branch_10__valid__0__anchor__out,
	output forkC_27__cst_7__valid__0__anchor__out,
	output [31 : 0] cst_2__icmp_9__data__0__anchor__out,
	output forkC_27__brCst_block6__data__0__anchor__out,
	output cst_2__icmp_9__ready__0__anchor__out,
	output phi_n11__branch_17__valid__0__anchor__out,
	output fork_8__store_0__valid__0__anchor__out,
	output branch_8__phi_n14__ready__0__anchor__out,
	output fork_18__branch_16__valid__0__anchor__out,
	output [31 : 0] fork_8__store_0__data__0__anchor__out,
	output fork_18__branch_18__valid__0__anchor__out,
	output fork_16__branch_8__ready__0__anchor__out,
	output phiC_18__forkC_24__data__0__anchor__out,
	output branch_3__sink_3__valid__0__anchor__out,
	output phi_n14__fork_10__valid__0__anchor__out,
	output [31 : 0] branch_7__phi_n13__data__0__anchor__out,
	output branchC_26__sink_15__data__0__anchor__out,
	output phiC_20__branchC_25__valid__0__anchor__out,
	output [31 : 0] fork_4__branch_20__data__0__anchor__out,
	output phiC_17__forkC_23__data__0__anchor__out,
	output source_1__cst_2__valid__0__anchor__out,
	output MC_A__load_20__ready__0__anchor__out,
	output branch_8__phi_n14__valid__0__anchor__out,
	output cst_8__MC_A__ready__0__anchor__out,
	output [30 : 0] phi_n15__branch_13__data__0__anchor__out,
	output branchC_25__phiC_22__valid__0__anchor__out,
	output [30 : 0] fork_3__branch_19__data__0__anchor__out,
	output branchC_25__phiC_21__ready__0__anchor__out,
	output forkC_27__branchC_26__data__0__anchor__out,
	output phi_n15__branch_13__ready__0__anchor__out,
	output fork_19__branch_20__data__0__anchor__out,
	output branch_15__sink_7__valid__0__anchor__out,
	output fork_15__branch_6__valid__0__anchor__out,
	output fork_10__branch_12__valid__0__anchor__out,
	output icmp_0__fork_22__data__0__anchor__out,
	output branch_18__Buffer_53__ready__0__anchor__out,
	output cst_0__icmp_0__valid__0__anchor__out,
	output [31 : 0] load_6__MC_A__data__0__anchor__out,
	output [31 : 0] phi_n16__branch_14__data__0__anchor__out,
	output cst_7__MC_A__valid__0__anchor__out,
	output fork_0__icmp_0__valid__0__anchor__out,
	output [31 : 0] branch_0__sink_0__data__0__anchor__out,
	output [31 : 0] Buffer_53__phi_n8__data__0__anchor__out,
	output forkC_24__branchC_23__data__0__anchor__out,
	output [31 : 0] load_20__MC_A__data__0__anchor__out,
	output [31 : 0] branch_15__sink_7__data__0__anchor__out,
	output forkC_24__branchC_23__valid__0__anchor__out,
	output branch_19__Buffer_52__ready__0__anchor__out,
	output end_valid,
	output fork_10__branch_12__ready__0__anchor__out,
	output phi_n9__fork_8__valid__0__anchor__out,
	output phi_n12__branch_18__valid__0__anchor__out,
	output load_14__MC_A__ready__0__anchor__out,
	output fork_18__branch_18__ready__0__anchor__out,
	output [31 : 0] A_dout0,
	output store_1__MC_A__valid__1__anchor__out,
	output branch_20__Buffer_50__ready__0__anchor__out,
	output branchC_21__phiC_17__ready__0__anchor__out,
	output phi_n5__fork_4__valid__0__anchor__out,
	output branch_4__sink_4__valid__0__anchor__out,
	output branchC_22__sink_13__ready__0__anchor__out,
	output brCst_block6__fork_18__data__0__anchor__out,
	output start_0__branchC_21__ready__0__anchor__out,
	output branchC_23__sink_14__data__0__anchor__out,
	output fork_17__branch_14__data__0__anchor__out,
	output [30 : 0] Buffer_52__phi_3__data__0__anchor__out,
	output [31 : 0] branch_14__phi_n5__data__0__anchor__out,
	output phiC_17__forkC_23__valid__0__anchor__out,
	output [30 : 0] add_27__fork_3__data__0__anchor__out,
	output [30 : 0] phi_n4__add_27__data__0__anchor__out,
	output phiC_19__phi_8__ready__0__anchor__out,
	output [31 : 0] branch_18__Buffer_53__data__0__anchor__out,
	output branch_4__phi_n8__valid__0__anchor__out,
	output cst_8__MC_A__valid__0__anchor__out,
	output MC_A__load_6__valid__0__anchor__out,
	output forkC_23__cst_1__data__0__anchor__out,
	output MC_A__end_0__data__0__anchor__out,
	output branch_9__phi_n15__valid__0__anchor__out,
	output fork_18__branchC_26__valid__0__anchor__out,
	output fork_14__branch_1__valid__0__anchor__out,
	output phiC_19__branchC_24__data__0__anchor__out,
	output cst_5__add_23__ready__0__anchor__out,
	output branch_1__sink_1__ready__0__anchor__out,
	output branch_19__sink_11__valid__0__anchor__out,
	output [31 : 0] MC_A__load_20__data__0__anchor__out,
	output source_1__cst_2__ready__0__anchor__out,
	output [31 : 0] phi_n10__branch_16__data__0__anchor__out,
	output cst_3__add_11__ready__0__anchor__out,
	output [31 : 0] A_dout1,
	output Buffer_56__phiC_18__ready__0__anchor__out,
	output [31 : 0] store_1__MC_A__data__0__anchor__out,
	output fork_2__branch_7__ready__0__anchor__out,
	output [31 : 0] fork_10__icmp_15__data__0__anchor__out,
	output fork_15__branchC_23__data__0__anchor__out,
	output icmp_28__fork_19__ready__0__anchor__out,
	output [31 : 0] n__fork_0__data__0__anchor__out,
	output fork_16__branchC_24__valid__0__anchor__out,
	output branch_16__sink_8__ready__0__anchor__out,
	output [31 : 0] phi_n13__fork_9__data__0__anchor__out,
	output fork_14__branchC_22__ready__0__anchor__out,
	output branch_5__sink_5__valid__0__anchor__out,
	output [31 : 0] store_0__MC_A__data__0__anchor__out,
	output forkC_27__cst_7__data__0__anchor__out,
	output fork_17__branch_13__data__0__anchor__out,
	output fork_17__branch_12__valid__0__anchor__out,
	output n_ready_in,
	output phiC_23__ret_0__ready__0__anchor__out,
	output [30 : 0] fork_1__branch_6__data__0__anchor__out,
	output fork_17__branch_13__valid__0__anchor__out,
	output phi_n7__branch_9__valid__0__anchor__out,
	output fork_17__branch_11__valid__0__anchor__out,
	output forkC_28__branchC_27__valid__0__anchor__out,
	output branch_6__sink_6__valid__0__anchor__out,
	output phi_n14__fork_10__ready__0__anchor__out,
	output forkC_23__branchC_22__data__0__anchor__out,
	output [31 : 0] store_1__MC_A__data__1__anchor__out,
	output branchC_24__phiC_20__ready__0__anchor__out,
	output branch_7__phi_n3__ready__0__anchor__out,
	output [31 : 0] branch_14__phi_n12__data__0__anchor__out,
	output phi_n11__branch_17__ready__0__anchor__out,
	output fork_22__branch_0__ready__0__anchor__out,
	output fork_15__branchC_23__valid__0__anchor__out,
	output fork_1__branch_6__valid__0__anchor__out,
	output [31 : 0] fork_3__icmp_28__data__0__anchor__out,
	output cst_5__add_23__valid__0__anchor__out,
	output [30 : 0] branch_9__phi_n15__data__0__anchor__out,
	output Buffer_53__phi_n8__ready__0__anchor__out,
	output brCst_block2__fork_14__valid__0__anchor__out,
	output A_we1,
	output phi_n16__branch_14__valid__0__anchor__out,
	output branch_17__Buffer_54__valid__0__anchor__out,
	output fork_9__branch_11__ready__0__anchor__out,
	output fork_17__branch_12__data__0__anchor__out,
	output branch_3__phi_n6__valid__0__anchor__out,
	output branch_5__phi_n7__valid__0__anchor__out,
	output [31 : 0] branch_16__Buffer_55__data__0__anchor__out,
	output store_1__MC_A__ready__0__anchor__out,
	output fork_15__branch_3__data__0__anchor__out,
	output phiC_21__forkC_27__data__0__anchor__out,
	output branch_20__sink_12__valid__0__anchor__out,
	output branch_16__Buffer_55__valid__0__anchor__out,
	output [30 : 0] cst_6__add_27__data__0__anchor__out,
	output branchC_24__phiC_22__data__0__anchor__out,
	output add_23__branch_15__ready__0__anchor__out,
	output icmp_15__Buffer_58__valid__0__anchor__out,
	output store_0__MC_A__valid__1__anchor__out,
	output source_2__cst_3__ready__0__anchor__out,
	output forkC_24__brCst_block3__ready__0__anchor__out,
	output fork_18__branch_16__data__0__anchor__out,
	output [30 : 0] fork_1__branch_5__data__0__anchor__out,
	output phi_n8__branch_10__ready__0__anchor__out,
	output [31 : 0] phi_n2__store_1__data__0__anchor__out,
	output fork_9__add_11__ready__0__anchor__out,
	output fork_1__load_6__valid__0__anchor__out,
	output fork_3__branch_19__valid__0__anchor__out,
	output Buffer_54__phi_n7__valid__0__anchor__out,
	output brCst_block6__fork_18__ready__0__anchor__out
);
	wire Buffer_58_clk;
	wire Buffer_58_rst;
	wire [31 : 0] Buffer_58_in1_data;
	wire Buffer_58_in1_ready;
	wire Buffer_58_in1_valid;
	wire [31 : 0] Buffer_58_out1_data;
	wire Buffer_58_out1_ready;
	wire Buffer_58_out1_valid;
	wire n_clk;
	wire n_rst;
	wire [31 : 0] n_in1_data;
	wire n_in1_ready;
	wire n_in1_valid;
	wire [31 : 0] n_out1_data;
	wire n_out1_ready;
	wire n_out1_valid;
	wire cst_0_clk;
	wire cst_0_rst;
	wire [1 : 0] cst_0_in1_data;
	wire cst_0_in1_ready;
	wire cst_0_in1_valid;
	wire [1 : 0] cst_0_out1_data;
	wire cst_0_out1_ready;
	wire cst_0_out1_valid;
	wire icmp_0_clk;
	wire icmp_0_rst;
	wire [31 : 0] icmp_0_in1_data;
	wire icmp_0_in1_ready;
	wire icmp_0_in1_valid;
	wire [31 : 0] icmp_0_in2_data;
	wire icmp_0_in2_ready;
	wire icmp_0_in2_valid;
	wire icmp_0_out1_data;
	wire icmp_0_out1_ready;
	wire icmp_0_out1_valid;
	wire brCst_block2_clk;
	wire brCst_block2_rst;
	wire brCst_block2_in1_data;
	wire brCst_block2_in1_ready;
	wire brCst_block2_in1_valid;
	wire brCst_block2_out1_data;
	wire brCst_block2_out1_ready;
	wire brCst_block2_out1_valid;
	wire cst_1_clk;
	wire cst_1_rst;
	wire cst_1_in1_data;
	wire cst_1_in1_ready;
	wire cst_1_in1_valid;
	wire cst_1_out1_data;
	wire cst_1_out1_ready;
	wire cst_1_out1_valid;
	wire phi_3_clk;
	wire phi_3_rst;
	wire phi_3_in1_data;
	wire phi_3_in1_ready;
	wire phi_3_in1_valid;
	wire [30 : 0] phi_3_in2_data;
	wire phi_3_in2_ready;
	wire phi_3_in2_valid;
	wire [30 : 0] phi_3_in3_data;
	wire phi_3_in3_ready;
	wire phi_3_in3_valid;
	wire [30 : 0] phi_3_out1_data;
	wire phi_3_out1_ready;
	wire phi_3_out1_valid;
	wire load_6_clk;
	wire load_6_rst;
	wire [31 : 0] load_6_in1_data;
	wire load_6_in1_ready;
	wire load_6_in1_valid;
	wire [30 : 0] load_6_in2_data;
	wire load_6_in2_ready;
	wire load_6_in2_valid;
	wire [31 : 0] load_6_out1_data;
	wire load_6_out1_ready;
	wire load_6_out1_valid;
	wire [30 : 0] load_6_out2_data;
	wire load_6_out2_ready;
	wire load_6_out2_valid;
	wire brCst_block3_clk;
	wire brCst_block3_rst;
	wire brCst_block3_in1_data;
	wire brCst_block3_in1_ready;
	wire brCst_block3_in1_valid;
	wire brCst_block3_out1_data;
	wire brCst_block3_out1_ready;
	wire brCst_block3_out1_valid;
	wire phi_8_clk;
	wire phi_8_rst;
	wire phi_8_in1_data;
	wire phi_8_in1_ready;
	wire phi_8_in1_valid;
	wire [31 : 0] phi_8_in2_data;
	wire phi_8_in2_ready;
	wire phi_8_in2_valid;
	wire [31 : 0] phi_8_in3_data;
	wire phi_8_in3_ready;
	wire phi_8_in3_valid;
	wire [31 : 0] phi_8_out1_data;
	wire phi_8_out1_ready;
	wire phi_8_out1_valid;
	wire cst_2_clk;
	wire cst_2_rst;
	wire cst_2_in1_data;
	wire cst_2_in1_ready;
	wire cst_2_in1_valid;
	wire cst_2_out1_data;
	wire cst_2_out1_ready;
	wire cst_2_out1_valid;
	wire icmp_9_clk;
	wire icmp_9_rst;
	wire [31 : 0] icmp_9_in1_data;
	wire icmp_9_in1_ready;
	wire icmp_9_in1_valid;
	wire [31 : 0] icmp_9_in2_data;
	wire icmp_9_in2_ready;
	wire icmp_9_in2_valid;
	wire icmp_9_out1_data;
	wire icmp_9_out1_ready;
	wire icmp_9_out1_valid;
	wire cst_3_clk;
	wire cst_3_rst;
	wire [31 : 0] cst_3_in1_data;
	wire cst_3_in1_ready;
	wire cst_3_in1_valid;
	wire [31 : 0] cst_3_out1_data;
	wire cst_3_out1_ready;
	wire cst_3_out1_valid;
	wire add_11_clk;
	wire add_11_rst;
	wire [31 : 0] add_11_in1_data;
	wire add_11_in1_ready;
	wire add_11_in1_valid;
	wire [31 : 0] add_11_in2_data;
	wire add_11_in2_ready;
	wire add_11_in2_valid;
	wire [31 : 0] add_11_out1_data;
	wire add_11_out1_ready;
	wire add_11_out1_valid;
	wire load_14_clk;
	wire load_14_rst;
	wire [31 : 0] load_14_in1_data;
	wire load_14_in1_ready;
	wire load_14_in1_valid;
	wire [31 : 0] load_14_in2_data;
	wire load_14_in2_ready;
	wire load_14_in2_valid;
	wire [31 : 0] load_14_out1_data;
	wire load_14_out1_ready;
	wire load_14_out1_valid;
	wire [31 : 0] load_14_out2_data;
	wire load_14_out2_ready;
	wire load_14_out2_valid;
	wire icmp_15_clk;
	wire icmp_15_rst;
	wire [31 : 0] icmp_15_in1_data;
	wire icmp_15_in1_ready;
	wire icmp_15_in1_valid;
	wire [31 : 0] icmp_15_in2_data;
	wire icmp_15_in2_ready;
	wire icmp_15_in2_valid;
	wire icmp_15_out1_data;
	wire icmp_15_out1_ready;
	wire icmp_15_out1_valid;
	wire cst_4_clk;
	wire cst_4_rst;
	wire [31 : 0] cst_4_in1_data;
	wire cst_4_in1_ready;
	wire cst_4_in1_valid;
	wire [31 : 0] cst_4_out1_data;
	wire cst_4_out1_ready;
	wire cst_4_out1_valid;
	wire add_17_clk;
	wire add_17_rst;
	wire [31 : 0] add_17_in1_data;
	wire add_17_in1_ready;
	wire add_17_in1_valid;
	wire [31 : 0] add_17_in2_data;
	wire add_17_in2_ready;
	wire add_17_in2_valid;
	wire [31 : 0] add_17_out1_data;
	wire add_17_out1_ready;
	wire add_17_out1_valid;
	wire load_20_clk;
	wire load_20_rst;
	wire [31 : 0] load_20_in1_data;
	wire load_20_in1_ready;
	wire load_20_in1_valid;
	wire [31 : 0] load_20_in2_data;
	wire load_20_in2_ready;
	wire load_20_in2_valid;
	wire [31 : 0] load_20_out1_data;
	wire load_20_out1_ready;
	wire load_20_out1_valid;
	wire [31 : 0] load_20_out2_data;
	wire load_20_out2_ready;
	wire load_20_out2_valid;
	wire store_0_clk;
	wire store_0_rst;
	wire [31 : 0] store_0_in1_data;
	wire store_0_in1_ready;
	wire store_0_in1_valid;
	wire [31 : 0] store_0_in2_data;
	wire store_0_in2_ready;
	wire store_0_in2_valid;
	wire [31 : 0] store_0_out1_data;
	wire store_0_out1_ready;
	wire store_0_out1_valid;
	wire [31 : 0] store_0_out2_data;
	wire store_0_out2_ready;
	wire store_0_out2_valid;
	wire cst_5_clk;
	wire cst_5_rst;
	wire [31 : 0] cst_5_in1_data;
	wire cst_5_in1_ready;
	wire cst_5_in1_valid;
	wire [31 : 0] cst_5_out1_data;
	wire cst_5_out1_ready;
	wire cst_5_out1_valid;
	wire add_23_clk;
	wire add_23_rst;
	wire [31 : 0] add_23_in1_data;
	wire add_23_in1_ready;
	wire add_23_in1_valid;
	wire [31 : 0] add_23_in2_data;
	wire add_23_in2_ready;
	wire add_23_in2_valid;
	wire [31 : 0] add_23_out1_data;
	wire add_23_out1_ready;
	wire add_23_out1_valid;
	wire brCst_block6_clk;
	wire brCst_block6_rst;
	wire brCst_block6_in1_data;
	wire brCst_block6_in1_ready;
	wire brCst_block6_in1_valid;
	wire brCst_block6_out1_data;
	wire brCst_block6_out1_ready;
	wire brCst_block6_out1_valid;
	wire store_1_clk;
	wire store_1_rst;
	wire [31 : 0] store_1_in1_data;
	wire store_1_in1_ready;
	wire store_1_in1_valid;
	wire [31 : 0] store_1_in2_data;
	wire store_1_in2_ready;
	wire store_1_in2_valid;
	wire [31 : 0] store_1_out1_data;
	wire store_1_out1_ready;
	wire store_1_out1_valid;
	wire [31 : 0] store_1_out2_data;
	wire store_1_out2_ready;
	wire store_1_out2_valid;
	wire cst_6_clk;
	wire cst_6_rst;
	wire cst_6_in1_data;
	wire cst_6_in1_ready;
	wire cst_6_in1_valid;
	wire cst_6_out1_data;
	wire cst_6_out1_ready;
	wire cst_6_out1_valid;
	wire add_27_clk;
	wire add_27_rst;
	wire [30 : 0] add_27_in1_data;
	wire add_27_in1_ready;
	wire add_27_in1_valid;
	wire [30 : 0] add_27_in2_data;
	wire add_27_in2_ready;
	wire add_27_in2_valid;
	wire [30 : 0] add_27_out1_data;
	wire add_27_out1_ready;
	wire add_27_out1_valid;
	wire icmp_28_clk;
	wire icmp_28_rst;
	wire [31 : 0] icmp_28_in1_data;
	wire icmp_28_in1_ready;
	wire icmp_28_in1_valid;
	wire [31 : 0] icmp_28_in2_data;
	wire icmp_28_in2_ready;
	wire icmp_28_in2_valid;
	wire icmp_28_out1_data;
	wire icmp_28_out1_ready;
	wire icmp_28_out1_valid;
	wire ret_0_clk;
	wire ret_0_rst;
	wire ret_0_in1_data;
	wire ret_0_in1_ready;
	wire ret_0_in1_valid;
	wire ret_0_out1_data;
	wire ret_0_out1_ready;
	wire ret_0_out1_valid;
	wire phi_n0_clk;
	wire phi_n0_rst;
	wire [31 : 0] phi_n0_in1_data;
	wire phi_n0_in1_ready;
	wire phi_n0_in1_valid;
	wire [31 : 0] phi_n0_out1_data;
	wire phi_n0_out1_ready;
	wire phi_n0_out1_valid;
	wire phi_n1_clk;
	wire phi_n1_rst;
	wire [31 : 0] phi_n1_in1_data;
	wire phi_n1_in1_ready;
	wire phi_n1_in1_valid;
	wire [31 : 0] phi_n1_in2_data;
	wire phi_n1_in2_ready;
	wire phi_n1_in2_valid;
	wire [31 : 0] phi_n1_out1_data;
	wire phi_n1_out1_ready;
	wire phi_n1_out1_valid;
	wire phi_n2_clk;
	wire phi_n2_rst;
	wire [31 : 0] phi_n2_in1_data;
	wire phi_n2_in1_ready;
	wire phi_n2_in1_valid;
	wire [31 : 0] phi_n2_in2_data;
	wire phi_n2_in2_ready;
	wire phi_n2_in2_valid;
	wire [31 : 0] phi_n2_out1_data;
	wire phi_n2_out1_ready;
	wire phi_n2_out1_valid;
	wire phi_n3_clk;
	wire phi_n3_rst;
	wire [31 : 0] phi_n3_in1_data;
	wire phi_n3_in1_ready;
	wire phi_n3_in1_valid;
	wire [31 : 0] phi_n3_in2_data;
	wire phi_n3_in2_ready;
	wire phi_n3_in2_valid;
	wire [31 : 0] phi_n3_out1_data;
	wire phi_n3_out1_ready;
	wire phi_n3_out1_valid;
	wire phi_n4_clk;
	wire phi_n4_rst;
	wire [30 : 0] phi_n4_in1_data;
	wire phi_n4_in1_ready;
	wire phi_n4_in1_valid;
	wire [30 : 0] phi_n4_in2_data;
	wire phi_n4_in2_ready;
	wire phi_n4_in2_valid;
	wire [30 : 0] phi_n4_out1_data;
	wire phi_n4_out1_ready;
	wire phi_n4_out1_valid;
	wire phi_n5_clk;
	wire phi_n5_rst;
	wire [31 : 0] phi_n5_in1_data;
	wire phi_n5_in1_ready;
	wire phi_n5_in1_valid;
	wire [31 : 0] phi_n5_in2_data;
	wire phi_n5_in2_ready;
	wire phi_n5_in2_valid;
	wire [31 : 0] phi_n5_out1_data;
	wire phi_n5_out1_ready;
	wire phi_n5_out1_valid;
	wire phi_n6_clk;
	wire phi_n6_rst;
	wire [31 : 0] phi_n6_in1_data;
	wire phi_n6_in1_ready;
	wire phi_n6_in1_valid;
	wire [31 : 0] phi_n6_in2_data;
	wire phi_n6_in2_ready;
	wire phi_n6_in2_valid;
	wire [31 : 0] phi_n6_out1_data;
	wire phi_n6_out1_ready;
	wire phi_n6_out1_valid;
	wire phi_n7_clk;
	wire phi_n7_rst;
	wire [30 : 0] phi_n7_in1_data;
	wire phi_n7_in1_ready;
	wire phi_n7_in1_valid;
	wire [30 : 0] phi_n7_in2_data;
	wire phi_n7_in2_ready;
	wire phi_n7_in2_valid;
	wire [30 : 0] phi_n7_out1_data;
	wire phi_n7_out1_ready;
	wire phi_n7_out1_valid;
	wire phi_n8_clk;
	wire phi_n8_rst;
	wire [31 : 0] phi_n8_in1_data;
	wire phi_n8_in1_ready;
	wire phi_n8_in1_valid;
	wire [31 : 0] phi_n8_in2_data;
	wire phi_n8_in2_ready;
	wire phi_n8_in2_valid;
	wire [31 : 0] phi_n8_out1_data;
	wire phi_n8_out1_ready;
	wire phi_n8_out1_valid;
	wire phi_n9_clk;
	wire phi_n9_rst;
	wire [31 : 0] phi_n9_in1_data;
	wire phi_n9_in1_ready;
	wire phi_n9_in1_valid;
	wire [31 : 0] phi_n9_out1_data;
	wire phi_n9_out1_ready;
	wire phi_n9_out1_valid;
	wire phi_n10_clk;
	wire phi_n10_rst;
	wire [31 : 0] phi_n10_in1_data;
	wire phi_n10_in1_ready;
	wire phi_n10_in1_valid;
	wire [31 : 0] phi_n10_out1_data;
	wire phi_n10_out1_ready;
	wire phi_n10_out1_valid;
	wire phi_n11_clk;
	wire phi_n11_rst;
	wire [30 : 0] phi_n11_in1_data;
	wire phi_n11_in1_ready;
	wire phi_n11_in1_valid;
	wire [30 : 0] phi_n11_out1_data;
	wire phi_n11_out1_ready;
	wire phi_n11_out1_valid;
	wire phi_n12_clk;
	wire phi_n12_rst;
	wire [31 : 0] phi_n12_in1_data;
	wire phi_n12_in1_ready;
	wire phi_n12_in1_valid;
	wire [31 : 0] phi_n12_out1_data;
	wire phi_n12_out1_ready;
	wire phi_n12_out1_valid;
	wire phi_n13_clk;
	wire phi_n13_rst;
	wire [31 : 0] phi_n13_in1_data;
	wire phi_n13_in1_ready;
	wire phi_n13_in1_valid;
	wire [31 : 0] phi_n13_out1_data;
	wire phi_n13_out1_ready;
	wire phi_n13_out1_valid;
	wire phi_n14_clk;
	wire phi_n14_rst;
	wire [31 : 0] phi_n14_in1_data;
	wire phi_n14_in1_ready;
	wire phi_n14_in1_valid;
	wire [31 : 0] phi_n14_out1_data;
	wire phi_n14_out1_ready;
	wire phi_n14_out1_valid;
	wire phi_n15_clk;
	wire phi_n15_rst;
	wire [30 : 0] phi_n15_in1_data;
	wire phi_n15_in1_ready;
	wire phi_n15_in1_valid;
	wire [30 : 0] phi_n15_out1_data;
	wire phi_n15_out1_ready;
	wire phi_n15_out1_valid;
	wire phi_n16_clk;
	wire phi_n16_rst;
	wire [31 : 0] phi_n16_in1_data;
	wire phi_n16_in1_ready;
	wire phi_n16_in1_valid;
	wire [31 : 0] phi_n16_out1_data;
	wire phi_n16_out1_ready;
	wire phi_n16_out1_valid;
	wire fork_0_clk;
	wire fork_0_rst;
	wire [31 : 0] fork_0_in1_data;
	wire fork_0_in1_ready;
	wire fork_0_in1_valid;
	wire [31 : 0] fork_0_out1_data;
	wire fork_0_out1_ready;
	wire fork_0_out1_valid;
	wire [31 : 0] fork_0_out2_data;
	wire fork_0_out2_ready;
	wire fork_0_out2_valid;
	wire fork_1_clk;
	wire fork_1_rst;
	wire [30 : 0] fork_1_in1_data;
	wire fork_1_in1_ready;
	wire fork_1_in1_valid;
	wire [30 : 0] fork_1_out1_data;
	wire fork_1_out1_ready;
	wire fork_1_out1_valid;
	wire [30 : 0] fork_1_out2_data;
	wire fork_1_out2_ready;
	wire fork_1_out2_valid;
	wire [30 : 0] fork_1_out3_data;
	wire fork_1_out3_ready;
	wire fork_1_out3_valid;
	wire fork_2_clk;
	wire fork_2_rst;
	wire [31 : 0] fork_2_in1_data;
	wire fork_2_in1_ready;
	wire fork_2_in1_valid;
	wire [31 : 0] fork_2_out1_data;
	wire fork_2_out1_ready;
	wire fork_2_out1_valid;
	wire [31 : 0] fork_2_out2_data;
	wire fork_2_out2_ready;
	wire fork_2_out2_valid;
	wire fork_3_clk;
	wire fork_3_rst;
	wire [30 : 0] fork_3_in1_data;
	wire fork_3_in1_ready;
	wire fork_3_in1_valid;
	wire [30 : 0] fork_3_out1_data;
	wire fork_3_out1_ready;
	wire fork_3_out1_valid;
	wire [30 : 0] fork_3_out2_data;
	wire fork_3_out2_ready;
	wire fork_3_out2_valid;
	wire fork_4_clk;
	wire fork_4_rst;
	wire [31 : 0] fork_4_in1_data;
	wire fork_4_in1_ready;
	wire fork_4_in1_valid;
	wire [31 : 0] fork_4_out1_data;
	wire fork_4_out1_ready;
	wire fork_4_out1_valid;
	wire [31 : 0] fork_4_out2_data;
	wire fork_4_out2_ready;
	wire fork_4_out2_valid;
	wire fork_8_clk;
	wire fork_8_rst;
	wire [31 : 0] fork_8_in1_data;
	wire fork_8_in1_ready;
	wire fork_8_in1_valid;
	wire [31 : 0] fork_8_out1_data;
	wire fork_8_out1_ready;
	wire fork_8_out1_valid;
	wire [31 : 0] fork_8_out2_data;
	wire fork_8_out2_ready;
	wire fork_8_out2_valid;
	wire [31 : 0] fork_8_out3_data;
	wire fork_8_out3_ready;
	wire fork_8_out3_valid;
	wire fork_9_clk;
	wire fork_9_rst;
	wire [31 : 0] fork_9_in1_data;
	wire fork_9_in1_ready;
	wire fork_9_in1_valid;
	wire [31 : 0] fork_9_out1_data;
	wire fork_9_out1_ready;
	wire fork_9_out1_valid;
	wire [31 : 0] fork_9_out2_data;
	wire fork_9_out2_ready;
	wire fork_9_out2_valid;
	wire fork_10_clk;
	wire fork_10_rst;
	wire [31 : 0] fork_10_in1_data;
	wire fork_10_in1_ready;
	wire fork_10_in1_valid;
	wire [31 : 0] fork_10_out1_data;
	wire fork_10_out1_ready;
	wire fork_10_out1_valid;
	wire [31 : 0] fork_10_out2_data;
	wire fork_10_out2_ready;
	wire fork_10_out2_valid;
	wire branch_0_clk;
	wire branch_0_rst;
	wire [31 : 0] branch_0_in1_data;
	wire branch_0_in1_ready;
	wire branch_0_in1_valid;
	wire branch_0_in2_data;
	wire branch_0_in2_ready;
	wire branch_0_in2_valid;
	wire [31 : 0] branch_0_out1_data;
	wire branch_0_out1_ready;
	wire branch_0_out1_valid;
	wire [31 : 0] branch_0_out2_data;
	wire branch_0_out2_ready;
	wire branch_0_out2_valid;
	wire branch_1_clk;
	wire branch_1_rst;
	wire branch_1_in1_data;
	wire branch_1_in1_ready;
	wire branch_1_in1_valid;
	wire branch_1_in2_data;
	wire branch_1_in2_ready;
	wire branch_1_in2_valid;
	wire branch_1_out1_data;
	wire branch_1_out1_ready;
	wire branch_1_out1_valid;
	wire branch_1_out2_data;
	wire branch_1_out2_ready;
	wire branch_1_out2_valid;
	wire branch_2_clk;
	wire branch_2_rst;
	wire [31 : 0] branch_2_in1_data;
	wire branch_2_in1_ready;
	wire branch_2_in1_valid;
	wire branch_2_in2_data;
	wire branch_2_in2_ready;
	wire branch_2_in2_valid;
	wire [31 : 0] branch_2_out1_data;
	wire branch_2_out1_ready;
	wire branch_2_out1_valid;
	wire [31 : 0] branch_2_out2_data;
	wire branch_2_out2_ready;
	wire branch_2_out2_valid;
	wire fork_14_clk;
	wire fork_14_rst;
	wire fork_14_in1_data;
	wire fork_14_in1_ready;
	wire fork_14_in1_valid;
	wire fork_14_out1_data;
	wire fork_14_out1_ready;
	wire fork_14_out1_valid;
	wire fork_14_out2_data;
	wire fork_14_out2_ready;
	wire fork_14_out2_valid;
	wire fork_14_out3_data;
	wire fork_14_out3_ready;
	wire fork_14_out3_valid;
	wire branch_3_clk;
	wire branch_3_rst;
	wire [31 : 0] branch_3_in1_data;
	wire branch_3_in1_ready;
	wire branch_3_in1_valid;
	wire branch_3_in2_data;
	wire branch_3_in2_ready;
	wire branch_3_in2_valid;
	wire [31 : 0] branch_3_out1_data;
	wire branch_3_out1_ready;
	wire branch_3_out1_valid;
	wire [31 : 0] branch_3_out2_data;
	wire branch_3_out2_ready;
	wire branch_3_out2_valid;
	wire branch_4_clk;
	wire branch_4_rst;
	wire [31 : 0] branch_4_in1_data;
	wire branch_4_in1_ready;
	wire branch_4_in1_valid;
	wire branch_4_in2_data;
	wire branch_4_in2_ready;
	wire branch_4_in2_valid;
	wire [31 : 0] branch_4_out1_data;
	wire branch_4_out1_ready;
	wire branch_4_out1_valid;
	wire [31 : 0] branch_4_out2_data;
	wire branch_4_out2_ready;
	wire branch_4_out2_valid;
	wire branch_5_clk;
	wire branch_5_rst;
	wire [30 : 0] branch_5_in1_data;
	wire branch_5_in1_ready;
	wire branch_5_in1_valid;
	wire branch_5_in2_data;
	wire branch_5_in2_ready;
	wire branch_5_in2_valid;
	wire [30 : 0] branch_5_out1_data;
	wire branch_5_out1_ready;
	wire branch_5_out1_valid;
	wire [30 : 0] branch_5_out2_data;
	wire branch_5_out2_ready;
	wire branch_5_out2_valid;
	wire branch_6_clk;
	wire branch_6_rst;
	wire [30 : 0] branch_6_in1_data;
	wire branch_6_in1_ready;
	wire branch_6_in1_valid;
	wire branch_6_in2_data;
	wire branch_6_in2_ready;
	wire branch_6_in2_valid;
	wire [30 : 0] branch_6_out1_data;
	wire branch_6_out1_ready;
	wire branch_6_out1_valid;
	wire [30 : 0] branch_6_out2_data;
	wire branch_6_out2_ready;
	wire branch_6_out2_valid;
	wire fork_15_clk;
	wire fork_15_rst;
	wire fork_15_in1_data;
	wire fork_15_in1_ready;
	wire fork_15_in1_valid;
	wire fork_15_out1_data;
	wire fork_15_out1_ready;
	wire fork_15_out1_valid;
	wire fork_15_out2_data;
	wire fork_15_out2_ready;
	wire fork_15_out2_valid;
	wire fork_15_out3_data;
	wire fork_15_out3_ready;
	wire fork_15_out3_valid;
	wire fork_15_out4_data;
	wire fork_15_out4_ready;
	wire fork_15_out4_valid;
	wire fork_15_out5_data;
	wire fork_15_out5_ready;
	wire fork_15_out5_valid;
	wire branch_7_clk;
	wire branch_7_rst;
	wire [31 : 0] branch_7_in1_data;
	wire branch_7_in1_ready;
	wire branch_7_in1_valid;
	wire branch_7_in2_data;
	wire branch_7_in2_ready;
	wire branch_7_in2_valid;
	wire [31 : 0] branch_7_out1_data;
	wire branch_7_out1_ready;
	wire branch_7_out1_valid;
	wire [31 : 0] branch_7_out2_data;
	wire branch_7_out2_ready;
	wire branch_7_out2_valid;
	wire branch_8_clk;
	wire branch_8_rst;
	wire [31 : 0] branch_8_in1_data;
	wire branch_8_in1_ready;
	wire branch_8_in1_valid;
	wire branch_8_in2_data;
	wire branch_8_in2_ready;
	wire branch_8_in2_valid;
	wire [31 : 0] branch_8_out1_data;
	wire branch_8_out1_ready;
	wire branch_8_out1_valid;
	wire [31 : 0] branch_8_out2_data;
	wire branch_8_out2_ready;
	wire branch_8_out2_valid;
	wire branch_9_clk;
	wire branch_9_rst;
	wire [30 : 0] branch_9_in1_data;
	wire branch_9_in1_ready;
	wire branch_9_in1_valid;
	wire branch_9_in2_data;
	wire branch_9_in2_ready;
	wire branch_9_in2_valid;
	wire [30 : 0] branch_9_out1_data;
	wire branch_9_out1_ready;
	wire branch_9_out1_valid;
	wire [30 : 0] branch_9_out2_data;
	wire branch_9_out2_ready;
	wire branch_9_out2_valid;
	wire branch_10_clk;
	wire branch_10_rst;
	wire [31 : 0] branch_10_in1_data;
	wire branch_10_in1_ready;
	wire branch_10_in1_valid;
	wire branch_10_in2_data;
	wire branch_10_in2_ready;
	wire branch_10_in2_valid;
	wire [31 : 0] branch_10_out1_data;
	wire branch_10_out1_ready;
	wire branch_10_out1_valid;
	wire [31 : 0] branch_10_out2_data;
	wire branch_10_out2_ready;
	wire branch_10_out2_valid;
	wire fork_16_clk;
	wire fork_16_rst;
	wire fork_16_in1_data;
	wire fork_16_in1_ready;
	wire fork_16_in1_valid;
	wire fork_16_out1_data;
	wire fork_16_out1_ready;
	wire fork_16_out1_valid;
	wire fork_16_out2_data;
	wire fork_16_out2_ready;
	wire fork_16_out2_valid;
	wire fork_16_out3_data;
	wire fork_16_out3_ready;
	wire fork_16_out3_valid;
	wire fork_16_out4_data;
	wire fork_16_out4_ready;
	wire fork_16_out4_valid;
	wire fork_16_out5_data;
	wire fork_16_out5_ready;
	wire fork_16_out5_valid;
	wire branch_11_clk;
	wire branch_11_rst;
	wire [31 : 0] branch_11_in1_data;
	wire branch_11_in1_ready;
	wire branch_11_in1_valid;
	wire branch_11_in2_data;
	wire branch_11_in2_ready;
	wire branch_11_in2_valid;
	wire [31 : 0] branch_11_out1_data;
	wire branch_11_out1_ready;
	wire branch_11_out1_valid;
	wire [31 : 0] branch_11_out2_data;
	wire branch_11_out2_ready;
	wire branch_11_out2_valid;
	wire branch_12_clk;
	wire branch_12_rst;
	wire [31 : 0] branch_12_in1_data;
	wire branch_12_in1_ready;
	wire branch_12_in1_valid;
	wire branch_12_in2_data;
	wire branch_12_in2_ready;
	wire branch_12_in2_valid;
	wire [31 : 0] branch_12_out1_data;
	wire branch_12_out1_ready;
	wire branch_12_out1_valid;
	wire [31 : 0] branch_12_out2_data;
	wire branch_12_out2_ready;
	wire branch_12_out2_valid;
	wire branch_13_clk;
	wire branch_13_rst;
	wire [30 : 0] branch_13_in1_data;
	wire branch_13_in1_ready;
	wire branch_13_in1_valid;
	wire branch_13_in2_data;
	wire branch_13_in2_ready;
	wire branch_13_in2_valid;
	wire [30 : 0] branch_13_out1_data;
	wire branch_13_out1_ready;
	wire branch_13_out1_valid;
	wire [30 : 0] branch_13_out2_data;
	wire branch_13_out2_ready;
	wire branch_13_out2_valid;
	wire branch_14_clk;
	wire branch_14_rst;
	wire [31 : 0] branch_14_in1_data;
	wire branch_14_in1_ready;
	wire branch_14_in1_valid;
	wire branch_14_in2_data;
	wire branch_14_in2_ready;
	wire branch_14_in2_valid;
	wire [31 : 0] branch_14_out1_data;
	wire branch_14_out1_ready;
	wire branch_14_out1_valid;
	wire [31 : 0] branch_14_out2_data;
	wire branch_14_out2_ready;
	wire branch_14_out2_valid;
	wire fork_17_clk;
	wire fork_17_rst;
	wire fork_17_in1_data;
	wire fork_17_in1_ready;
	wire fork_17_in1_valid;
	wire fork_17_out1_data;
	wire fork_17_out1_ready;
	wire fork_17_out1_valid;
	wire fork_17_out2_data;
	wire fork_17_out2_ready;
	wire fork_17_out2_valid;
	wire fork_17_out3_data;
	wire fork_17_out3_ready;
	wire fork_17_out3_valid;
	wire fork_17_out4_data;
	wire fork_17_out4_ready;
	wire fork_17_out4_valid;
	wire fork_17_out5_data;
	wire fork_17_out5_ready;
	wire fork_17_out5_valid;
	wire branch_15_clk;
	wire branch_15_rst;
	wire [31 : 0] branch_15_in1_data;
	wire branch_15_in1_ready;
	wire branch_15_in1_valid;
	wire branch_15_in2_data;
	wire branch_15_in2_ready;
	wire branch_15_in2_valid;
	wire [31 : 0] branch_15_out1_data;
	wire branch_15_out1_ready;
	wire branch_15_out1_valid;
	wire [31 : 0] branch_15_out2_data;
	wire branch_15_out2_ready;
	wire branch_15_out2_valid;
	wire branch_16_clk;
	wire branch_16_rst;
	wire [31 : 0] branch_16_in1_data;
	wire branch_16_in1_ready;
	wire branch_16_in1_valid;
	wire branch_16_in2_data;
	wire branch_16_in2_ready;
	wire branch_16_in2_valid;
	wire [31 : 0] branch_16_out1_data;
	wire branch_16_out1_ready;
	wire branch_16_out1_valid;
	wire [31 : 0] branch_16_out2_data;
	wire branch_16_out2_ready;
	wire branch_16_out2_valid;
	wire branch_17_clk;
	wire branch_17_rst;
	wire [30 : 0] branch_17_in1_data;
	wire branch_17_in1_ready;
	wire branch_17_in1_valid;
	wire branch_17_in2_data;
	wire branch_17_in2_ready;
	wire branch_17_in2_valid;
	wire [30 : 0] branch_17_out1_data;
	wire branch_17_out1_ready;
	wire branch_17_out1_valid;
	wire [30 : 0] branch_17_out2_data;
	wire branch_17_out2_ready;
	wire branch_17_out2_valid;
	wire branch_18_clk;
	wire branch_18_rst;
	wire [31 : 0] branch_18_in1_data;
	wire branch_18_in1_ready;
	wire branch_18_in1_valid;
	wire branch_18_in2_data;
	wire branch_18_in2_ready;
	wire branch_18_in2_valid;
	wire [31 : 0] branch_18_out1_data;
	wire branch_18_out1_ready;
	wire branch_18_out1_valid;
	wire [31 : 0] branch_18_out2_data;
	wire branch_18_out2_ready;
	wire branch_18_out2_valid;
	wire fork_18_clk;
	wire fork_18_rst;
	wire fork_18_in1_data;
	wire fork_18_in1_ready;
	wire fork_18_in1_valid;
	wire fork_18_out1_data;
	wire fork_18_out1_ready;
	wire fork_18_out1_valid;
	wire fork_18_out2_data;
	wire fork_18_out2_ready;
	wire fork_18_out2_valid;
	wire fork_18_out3_data;
	wire fork_18_out3_ready;
	wire fork_18_out3_valid;
	wire fork_18_out4_data;
	wire fork_18_out4_ready;
	wire fork_18_out4_valid;
	wire fork_18_out5_data;
	wire fork_18_out5_ready;
	wire fork_18_out5_valid;
	wire branch_19_clk;
	wire branch_19_rst;
	wire [30 : 0] branch_19_in1_data;
	wire branch_19_in1_ready;
	wire branch_19_in1_valid;
	wire branch_19_in2_data;
	wire branch_19_in2_ready;
	wire branch_19_in2_valid;
	wire [30 : 0] branch_19_out1_data;
	wire branch_19_out1_ready;
	wire branch_19_out1_valid;
	wire [30 : 0] branch_19_out2_data;
	wire branch_19_out2_ready;
	wire branch_19_out2_valid;
	wire branch_20_clk;
	wire branch_20_rst;
	wire [31 : 0] branch_20_in1_data;
	wire branch_20_in1_ready;
	wire branch_20_in1_valid;
	wire branch_20_in2_data;
	wire branch_20_in2_ready;
	wire branch_20_in2_valid;
	wire [31 : 0] branch_20_out1_data;
	wire branch_20_out1_ready;
	wire branch_20_out1_valid;
	wire [31 : 0] branch_20_out2_data;
	wire branch_20_out2_ready;
	wire branch_20_out2_valid;
	wire fork_19_clk;
	wire fork_19_rst;
	wire fork_19_in1_data;
	wire fork_19_in1_ready;
	wire fork_19_in1_valid;
	wire fork_19_out1_data;
	wire fork_19_out1_ready;
	wire fork_19_out1_valid;
	wire fork_19_out2_data;
	wire fork_19_out2_ready;
	wire fork_19_out2_valid;
	wire fork_19_out3_data;
	wire fork_19_out3_ready;
	wire fork_19_out3_valid;
	wire MC_A_clk;
	wire MC_A_rst;
	wire [31 : 0] MC_A_in1_data;
	wire MC_A_in1_ready;
	wire MC_A_in1_valid;
	wire [31 : 0] MC_A_in2_data;
	wire MC_A_in2_ready;
	wire MC_A_in2_valid;
	wire [31 : 0] MC_A_in3_data;
	wire MC_A_in3_ready;
	wire MC_A_in3_valid;
	wire [31 : 0] MC_A_in4_data;
	wire MC_A_in4_ready;
	wire MC_A_in4_valid;
	wire [31 : 0] MC_A_in5_data;
	wire MC_A_in5_ready;
	wire MC_A_in5_valid;
	wire [31 : 0] MC_A_in6_data;
	wire MC_A_in6_ready;
	wire MC_A_in6_valid;
	wire [31 : 0] MC_A_in7_data;
	wire MC_A_in7_ready;
	wire MC_A_in7_valid;
	wire [31 : 0] MC_A_in8_data;
	wire MC_A_in8_ready;
	wire MC_A_in8_valid;
	wire [31 : 0] MC_A_in9_data;
	wire MC_A_in9_ready;
	wire MC_A_in9_valid;
	wire [31 : 0] MC_A_out1_data;
	wire MC_A_out1_ready;
	wire MC_A_out1_valid;
	wire [31 : 0] MC_A_out2_data;
	wire MC_A_out2_ready;
	wire MC_A_out2_valid;
	wire [31 : 0] MC_A_out3_data;
	wire MC_A_out3_ready;
	wire MC_A_out3_valid;
	wire MC_A_out4_data;
	wire MC_A_out4_ready;
	wire MC_A_out4_valid;
	wire cst_7_clk;
	wire cst_7_rst;
	wire cst_7_in1_data;
	wire cst_7_in1_ready;
	wire cst_7_in1_valid;
	wire cst_7_out1_data;
	wire cst_7_out1_ready;
	wire cst_7_out1_valid;
	wire cst_8_clk;
	wire cst_8_rst;
	wire cst_8_in1_data;
	wire cst_8_in1_ready;
	wire cst_8_in1_valid;
	wire cst_8_out1_data;
	wire cst_8_out1_ready;
	wire cst_8_out1_valid;
	wire end_0_clk;
	wire end_0_rst;
	wire end_0_in1_data;
	wire end_0_in1_ready;
	wire end_0_in1_valid;
	wire end_0_in2_data;
	wire end_0_in2_ready;
	wire end_0_in2_valid;
	wire end_0_out1_data;
	wire end_0_out1_ready;
	wire end_0_out1_valid;
	wire start_0_clk;
	wire start_0_rst;
	wire start_0_in1_data;
	wire start_0_in1_ready;
	wire start_0_in1_valid;
	wire start_0_out1_data;
	wire start_0_out1_ready;
	wire start_0_out1_valid;
	wire branchC_21_clk;
	wire branchC_21_rst;
	wire branchC_21_in1_data;
	wire branchC_21_in1_ready;
	wire branchC_21_in1_valid;
	wire branchC_21_in2_data;
	wire branchC_21_in2_ready;
	wire branchC_21_in2_valid;
	wire branchC_21_out1_data;
	wire branchC_21_out1_ready;
	wire branchC_21_out1_valid;
	wire branchC_21_out2_data;
	wire branchC_21_out2_ready;
	wire branchC_21_out2_valid;
	wire fork_22_clk;
	wire fork_22_rst;
	wire fork_22_in1_data;
	wire fork_22_in1_ready;
	wire fork_22_in1_valid;
	wire fork_22_out1_data;
	wire fork_22_out1_ready;
	wire fork_22_out1_valid;
	wire fork_22_out2_data;
	wire fork_22_out2_ready;
	wire fork_22_out2_valid;
	wire phiC_17_clk;
	wire phiC_17_rst;
	wire phiC_17_in1_data;
	wire phiC_17_in1_ready;
	wire phiC_17_in1_valid;
	wire phiC_17_out1_data;
	wire phiC_17_out1_ready;
	wire phiC_17_out1_valid;
	wire forkC_23_clk;
	wire forkC_23_rst;
	wire forkC_23_in1_data;
	wire forkC_23_in1_ready;
	wire forkC_23_in1_valid;
	wire forkC_23_out1_data;
	wire forkC_23_out1_ready;
	wire forkC_23_out1_valid;
	wire forkC_23_out2_data;
	wire forkC_23_out2_ready;
	wire forkC_23_out2_valid;
	wire forkC_23_out3_data;
	wire forkC_23_out3_ready;
	wire forkC_23_out3_valid;
	wire branchC_22_clk;
	wire branchC_22_rst;
	wire branchC_22_in1_data;
	wire branchC_22_in1_ready;
	wire branchC_22_in1_valid;
	wire branchC_22_in2_data;
	wire branchC_22_in2_ready;
	wire branchC_22_in2_valid;
	wire branchC_22_out1_data;
	wire branchC_22_out1_ready;
	wire branchC_22_out1_valid;
	wire branchC_22_out2_data;
	wire branchC_22_out2_ready;
	wire branchC_22_out2_valid;
	wire phiC_18_clk;
	wire phiC_18_rst;
	wire phiC_18_in1_data;
	wire phiC_18_in1_ready;
	wire phiC_18_in1_valid;
	wire phiC_18_in2_data;
	wire phiC_18_in2_ready;
	wire phiC_18_in2_valid;
	wire phiC_18_out1_data;
	wire phiC_18_out1_ready;
	wire phiC_18_out1_valid;
	wire phiC_18_out2_data;
	wire phiC_18_out2_ready;
	wire phiC_18_out2_valid;
	wire forkC_24_clk;
	wire forkC_24_rst;
	wire forkC_24_in1_data;
	wire forkC_24_in1_ready;
	wire forkC_24_in1_valid;
	wire forkC_24_out1_data;
	wire forkC_24_out1_ready;
	wire forkC_24_out1_valid;
	wire forkC_24_out2_data;
	wire forkC_24_out2_ready;
	wire forkC_24_out2_valid;
	wire branchC_23_clk;
	wire branchC_23_rst;
	wire branchC_23_in1_data;
	wire branchC_23_in1_ready;
	wire branchC_23_in1_valid;
	wire branchC_23_in2_data;
	wire branchC_23_in2_ready;
	wire branchC_23_in2_valid;
	wire branchC_23_out1_data;
	wire branchC_23_out1_ready;
	wire branchC_23_out1_valid;
	wire branchC_23_out2_data;
	wire branchC_23_out2_ready;
	wire branchC_23_out2_valid;
	wire phiC_19_clk;
	wire phiC_19_rst;
	wire phiC_19_in1_data;
	wire phiC_19_in1_ready;
	wire phiC_19_in1_valid;
	wire phiC_19_in2_data;
	wire phiC_19_in2_ready;
	wire phiC_19_in2_valid;
	wire phiC_19_out1_data;
	wire phiC_19_out1_ready;
	wire phiC_19_out1_valid;
	wire phiC_19_out2_data;
	wire phiC_19_out2_ready;
	wire phiC_19_out2_valid;
	wire branchC_24_clk;
	wire branchC_24_rst;
	wire branchC_24_in1_data;
	wire branchC_24_in1_ready;
	wire branchC_24_in1_valid;
	wire branchC_24_in2_data;
	wire branchC_24_in2_ready;
	wire branchC_24_in2_valid;
	wire branchC_24_out1_data;
	wire branchC_24_out1_ready;
	wire branchC_24_out1_valid;
	wire branchC_24_out2_data;
	wire branchC_24_out2_ready;
	wire branchC_24_out2_valid;
	wire phiC_20_clk;
	wire phiC_20_rst;
	wire phiC_20_in1_data;
	wire phiC_20_in1_ready;
	wire phiC_20_in1_valid;
	wire phiC_20_out1_data;
	wire phiC_20_out1_ready;
	wire phiC_20_out1_valid;
	wire branchC_25_clk;
	wire branchC_25_rst;
	wire branchC_25_in1_data;
	wire branchC_25_in1_ready;
	wire branchC_25_in1_valid;
	wire branchC_25_in2_data;
	wire branchC_25_in2_ready;
	wire branchC_25_in2_valid;
	wire branchC_25_out1_data;
	wire branchC_25_out1_ready;
	wire branchC_25_out1_valid;
	wire branchC_25_out2_data;
	wire branchC_25_out2_ready;
	wire branchC_25_out2_valid;
	wire phiC_21_clk;
	wire phiC_21_rst;
	wire phiC_21_in1_data;
	wire phiC_21_in1_ready;
	wire phiC_21_in1_valid;
	wire phiC_21_out1_data;
	wire phiC_21_out1_ready;
	wire phiC_21_out1_valid;
	wire forkC_27_clk;
	wire forkC_27_rst;
	wire forkC_27_in1_data;
	wire forkC_27_in1_ready;
	wire forkC_27_in1_valid;
	wire forkC_27_out1_data;
	wire forkC_27_out1_ready;
	wire forkC_27_out1_valid;
	wire forkC_27_out2_data;
	wire forkC_27_out2_ready;
	wire forkC_27_out2_valid;
	wire forkC_27_out3_data;
	wire forkC_27_out3_ready;
	wire forkC_27_out3_valid;
	wire branchC_26_clk;
	wire branchC_26_rst;
	wire branchC_26_in1_data;
	wire branchC_26_in1_ready;
	wire branchC_26_in1_valid;
	wire branchC_26_in2_data;
	wire branchC_26_in2_ready;
	wire branchC_26_in2_valid;
	wire branchC_26_out1_data;
	wire branchC_26_out1_ready;
	wire branchC_26_out1_valid;
	wire branchC_26_out2_data;
	wire branchC_26_out2_ready;
	wire branchC_26_out2_valid;
	wire phiC_22_clk;
	wire phiC_22_rst;
	wire phiC_22_in1_data;
	wire phiC_22_in1_ready;
	wire phiC_22_in1_valid;
	wire phiC_22_in2_data;
	wire phiC_22_in2_ready;
	wire phiC_22_in2_valid;
	wire phiC_22_out1_data;
	wire phiC_22_out1_ready;
	wire phiC_22_out1_valid;
	wire forkC_28_clk;
	wire forkC_28_rst;
	wire forkC_28_in1_data;
	wire forkC_28_in1_ready;
	wire forkC_28_in1_valid;
	wire forkC_28_out1_data;
	wire forkC_28_out1_ready;
	wire forkC_28_out1_valid;
	wire forkC_28_out2_data;
	wire forkC_28_out2_ready;
	wire forkC_28_out2_valid;
	wire branchC_27_clk;
	wire branchC_27_rst;
	wire branchC_27_in1_data;
	wire branchC_27_in1_ready;
	wire branchC_27_in1_valid;
	wire branchC_27_in2_data;
	wire branchC_27_in2_ready;
	wire branchC_27_in2_valid;
	wire branchC_27_out1_data;
	wire branchC_27_out1_ready;
	wire branchC_27_out1_valid;
	wire branchC_27_out2_data;
	wire branchC_27_out2_ready;
	wire branchC_27_out2_valid;
	wire phiC_23_clk;
	wire phiC_23_rst;
	wire phiC_23_in1_data;
	wire phiC_23_in1_ready;
	wire phiC_23_in1_valid;
	wire phiC_23_in2_data;
	wire phiC_23_in2_ready;
	wire phiC_23_in2_valid;
	wire phiC_23_out1_data;
	wire phiC_23_out1_ready;
	wire phiC_23_out1_valid;
	wire sink_0_clk;
	wire sink_0_rst;
	wire [31 : 0] sink_0_in1_data;
	wire sink_0_in1_ready;
	wire sink_0_in1_valid;
	wire sink_1_clk;
	wire sink_1_rst;
	wire sink_1_in1_data;
	wire sink_1_in1_ready;
	wire sink_1_in1_valid;
	wire sink_2_clk;
	wire sink_2_rst;
	wire [31 : 0] sink_2_in1_data;
	wire sink_2_in1_ready;
	wire sink_2_in1_valid;
	wire sink_3_clk;
	wire sink_3_rst;
	wire [31 : 0] sink_3_in1_data;
	wire sink_3_in1_ready;
	wire sink_3_in1_valid;
	wire sink_4_clk;
	wire sink_4_rst;
	wire [31 : 0] sink_4_in1_data;
	wire sink_4_in1_ready;
	wire sink_4_in1_valid;
	wire sink_5_clk;
	wire sink_5_rst;
	wire [30 : 0] sink_5_in1_data;
	wire sink_5_in1_ready;
	wire sink_5_in1_valid;
	wire sink_6_clk;
	wire sink_6_rst;
	wire [30 : 0] sink_6_in1_data;
	wire sink_6_in1_ready;
	wire sink_6_in1_valid;
	wire sink_7_clk;
	wire sink_7_rst;
	wire [31 : 0] sink_7_in1_data;
	wire sink_7_in1_ready;
	wire sink_7_in1_valid;
	wire sink_8_clk;
	wire sink_8_rst;
	wire [31 : 0] sink_8_in1_data;
	wire sink_8_in1_ready;
	wire sink_8_in1_valid;
	wire sink_9_clk;
	wire sink_9_rst;
	wire [30 : 0] sink_9_in1_data;
	wire sink_9_in1_ready;
	wire sink_9_in1_valid;
	wire sink_10_clk;
	wire sink_10_rst;
	wire [31 : 0] sink_10_in1_data;
	wire sink_10_in1_ready;
	wire sink_10_in1_valid;
	wire sink_11_clk;
	wire sink_11_rst;
	wire [30 : 0] sink_11_in1_data;
	wire sink_11_in1_ready;
	wire sink_11_in1_valid;
	wire sink_12_clk;
	wire sink_12_rst;
	wire [31 : 0] sink_12_in1_data;
	wire sink_12_in1_ready;
	wire sink_12_in1_valid;
	wire sink_13_clk;
	wire sink_13_rst;
	wire sink_13_in1_data;
	wire sink_13_in1_ready;
	wire sink_13_in1_valid;
	wire sink_14_clk;
	wire sink_14_rst;
	wire sink_14_in1_data;
	wire sink_14_in1_ready;
	wire sink_14_in1_valid;
	wire sink_15_clk;
	wire sink_15_rst;
	wire sink_15_in1_data;
	wire sink_15_in1_ready;
	wire sink_15_in1_valid;
	wire source_0_clk;
	wire source_0_rst;
	wire [1 : 0] source_0_out1_data;
	wire source_0_out1_ready;
	wire source_0_out1_valid;
	wire source_1_clk;
	wire source_1_rst;
	wire source_1_out1_data;
	wire source_1_out1_ready;
	wire source_1_out1_valid;
	wire source_2_clk;
	wire source_2_rst;
	wire [31 : 0] source_2_out1_data;
	wire source_2_out1_ready;
	wire source_2_out1_valid;
	wire source_3_clk;
	wire source_3_rst;
	wire [31 : 0] source_3_out1_data;
	wire source_3_out1_ready;
	wire source_3_out1_valid;
	wire source_4_clk;
	wire source_4_rst;
	wire [31 : 0] source_4_out1_data;
	wire source_4_out1_ready;
	wire source_4_out1_valid;
	wire source_5_clk;
	wire source_5_rst;
	wire source_5_out1_data;
	wire source_5_out1_ready;
	wire source_5_out1_valid;
	wire Buffer_50_clk;
	wire Buffer_50_rst;
	wire [31 : 0] Buffer_50_in1_data;
	wire Buffer_50_in1_ready;
	wire Buffer_50_in1_valid;
	wire [31 : 0] Buffer_50_out1_data;
	wire Buffer_50_out1_ready;
	wire Buffer_50_out1_valid;
	wire Buffer_51_clk;
	wire Buffer_51_rst;
	wire [31 : 0] Buffer_51_in1_data;
	wire Buffer_51_in1_ready;
	wire Buffer_51_in1_valid;
	wire [31 : 0] Buffer_51_out1_data;
	wire Buffer_51_out1_ready;
	wire Buffer_51_out1_valid;
	wire Buffer_52_clk;
	wire Buffer_52_rst;
	wire [30 : 0] Buffer_52_in1_data;
	wire Buffer_52_in1_ready;
	wire Buffer_52_in1_valid;
	wire [30 : 0] Buffer_52_out1_data;
	wire Buffer_52_out1_ready;
	wire Buffer_52_out1_valid;
	wire Buffer_53_clk;
	wire Buffer_53_rst;
	wire [31 : 0] Buffer_53_in1_data;
	wire Buffer_53_in1_ready;
	wire Buffer_53_in1_valid;
	wire [31 : 0] Buffer_53_out1_data;
	wire Buffer_53_out1_ready;
	wire Buffer_53_out1_valid;
	wire Buffer_54_clk;
	wire Buffer_54_rst;
	wire [30 : 0] Buffer_54_in1_data;
	wire Buffer_54_in1_ready;
	wire Buffer_54_in1_valid;
	wire [30 : 0] Buffer_54_out1_data;
	wire Buffer_54_out1_ready;
	wire Buffer_54_out1_valid;
	wire Buffer_55_clk;
	wire Buffer_55_rst;
	wire [31 : 0] Buffer_55_in1_data;
	wire Buffer_55_in1_ready;
	wire Buffer_55_in1_valid;
	wire [31 : 0] Buffer_55_out1_data;
	wire Buffer_55_out1_ready;
	wire Buffer_55_out1_valid;
	wire Buffer_56_clk;
	wire Buffer_56_rst;
	wire Buffer_56_in1_data;
	wire Buffer_56_in1_ready;
	wire Buffer_56_in1_valid;
	wire Buffer_56_out1_data;
	wire Buffer_56_out1_ready;
	wire Buffer_56_out1_valid;
	wire Buffer_57_clk;
	wire Buffer_57_rst;
	wire Buffer_57_in1_data;
	wire Buffer_57_in1_ready;
	wire Buffer_57_in1_valid;
	wire Buffer_57_out1_data;
	wire Buffer_57_out1_ready;
	wire Buffer_57_out1_valid;
	assign Buffer_58_clk = clk;
	assign Buffer_58_rst = rst;
	assign fork_17_in1_data = Buffer_58__fork_17__data__0__anchor__in;
	assign Buffer_58__fork_17__data__0__anchor__out = Buffer_58_out1_data;
	assign fork_17_in1_valid = Buffer_58__fork_17__valid__0__anchor__in;
	assign Buffer_58__fork_17__valid__0__anchor__out = Buffer_58_out1_valid;
	assign Buffer_58_out1_ready = Buffer_58__fork_17__ready__0__anchor__in;
	assign Buffer_58__fork_17__ready__0__anchor__out = fork_17_in1_ready;
	assign n_clk = clk;
	assign n_rst = rst;
	assign n_in1_data = n_din;
	assign n_in1_valid = n_valid_in;
	assign n_ready_in = n_in1_ready;
	assign fork_0_in1_data = n__fork_0__data__0__anchor__in;
	assign n__fork_0__data__0__anchor__out = n_out1_data;
	assign fork_0_in1_valid = n__fork_0__valid__0__anchor__in;
	assign n__fork_0__valid__0__anchor__out = n_out1_valid;
	assign n_out1_ready = n__fork_0__ready__0__anchor__in;
	assign n__fork_0__ready__0__anchor__out = fork_0_in1_ready;
	assign cst_0_clk = clk;
	assign cst_0_rst = rst;
	assign icmp_0_in2_data = cst_0__icmp_0__data__0__anchor__in;
	assign cst_0__icmp_0__data__0__anchor__out = cst_0_out1_data;
	assign icmp_0_in2_valid = cst_0__icmp_0__valid__0__anchor__in;
	assign cst_0__icmp_0__valid__0__anchor__out = cst_0_out1_valid;
	assign cst_0_out1_ready = cst_0__icmp_0__ready__0__anchor__in;
	assign cst_0__icmp_0__ready__0__anchor__out = icmp_0_in2_ready;
	assign icmp_0_clk = clk;
	assign icmp_0_rst = rst;
	assign fork_22_in1_data = icmp_0__fork_22__data__0__anchor__in;
	assign icmp_0__fork_22__data__0__anchor__out = icmp_0_out1_data;
	assign fork_22_in1_valid = icmp_0__fork_22__valid__0__anchor__in;
	assign icmp_0__fork_22__valid__0__anchor__out = icmp_0_out1_valid;
	assign icmp_0_out1_ready = icmp_0__fork_22__ready__0__anchor__in;
	assign icmp_0__fork_22__ready__0__anchor__out = fork_22_in1_ready;
	assign brCst_block2_clk = clk;
	assign brCst_block2_rst = rst;
	assign fork_14_in1_data = brCst_block2__fork_14__data__0__anchor__in;
	assign brCst_block2__fork_14__data__0__anchor__out = brCst_block2_out1_data;
	assign fork_14_in1_valid = brCst_block2__fork_14__valid__0__anchor__in;
	assign brCst_block2__fork_14__valid__0__anchor__out = brCst_block2_out1_valid;
	assign brCst_block2_out1_ready = brCst_block2__fork_14__ready__0__anchor__in;
	assign brCst_block2__fork_14__ready__0__anchor__out = fork_14_in1_ready;
	assign cst_1_clk = clk;
	assign cst_1_rst = rst;
	assign branch_1_in1_data = cst_1__branch_1__data__0__anchor__in;
	assign cst_1__branch_1__data__0__anchor__out = cst_1_out1_data;
	assign branch_1_in1_valid = cst_1__branch_1__valid__0__anchor__in;
	assign cst_1__branch_1__valid__0__anchor__out = cst_1_out1_valid;
	assign cst_1_out1_ready = cst_1__branch_1__ready__0__anchor__in;
	assign cst_1__branch_1__ready__0__anchor__out = branch_1_in1_ready;
	assign phi_3_clk = clk;
	assign phi_3_rst = rst;
	assign fork_1_in1_data = phi_3__fork_1__data__0__anchor__in;
	assign phi_3__fork_1__data__0__anchor__out = phi_3_out1_data;
	assign fork_1_in1_valid = phi_3__fork_1__valid__0__anchor__in;
	assign phi_3__fork_1__valid__0__anchor__out = phi_3_out1_valid;
	assign phi_3_out1_ready = phi_3__fork_1__ready__0__anchor__in;
	assign phi_3__fork_1__ready__0__anchor__out = fork_1_in1_ready;
	assign load_6_clk = clk;
	assign load_6_rst = rst;
	assign branch_3_in1_data = load_6__branch_3__data__0__anchor__in;
	assign load_6__branch_3__data__0__anchor__out = load_6_out1_data;
	assign branch_3_in1_valid = load_6__branch_3__valid__0__anchor__in;
	assign load_6__branch_3__valid__0__anchor__out = load_6_out1_valid;
	assign load_6_out1_ready = load_6__branch_3__ready__0__anchor__in;
	assign load_6__branch_3__ready__0__anchor__out = branch_3_in1_ready;
	assign MC_A_in3_data = load_6__MC_A__data__0__anchor__in;
	assign load_6__MC_A__data__0__anchor__out = load_6_out2_data;
	assign MC_A_in3_valid = load_6__MC_A__valid__0__anchor__in;
	assign load_6__MC_A__valid__0__anchor__out = load_6_out2_valid;
	assign load_6_out2_ready = load_6__MC_A__ready__0__anchor__in;
	assign load_6__MC_A__ready__0__anchor__out = MC_A_in3_ready;
	assign brCst_block3_clk = clk;
	assign brCst_block3_rst = rst;
	assign fork_15_in1_data = brCst_block3__fork_15__data__0__anchor__in;
	assign brCst_block3__fork_15__data__0__anchor__out = brCst_block3_out1_data;
	assign fork_15_in1_valid = brCst_block3__fork_15__valid__0__anchor__in;
	assign brCst_block3__fork_15__valid__0__anchor__out = brCst_block3_out1_valid;
	assign brCst_block3_out1_ready = brCst_block3__fork_15__ready__0__anchor__in;
	assign brCst_block3__fork_15__ready__0__anchor__out = fork_15_in1_ready;
	assign phi_8_clk = clk;
	assign phi_8_rst = rst;
	assign fork_2_in1_data = phi_8__fork_2__data__0__anchor__in;
	assign phi_8__fork_2__data__0__anchor__out = phi_8_out1_data;
	assign fork_2_in1_valid = phi_8__fork_2__valid__0__anchor__in;
	assign phi_8__fork_2__valid__0__anchor__out = phi_8_out1_valid;
	assign phi_8_out1_ready = phi_8__fork_2__ready__0__anchor__in;
	assign phi_8__fork_2__ready__0__anchor__out = fork_2_in1_ready;
	assign cst_2_clk = clk;
	assign cst_2_rst = rst;
	assign icmp_9_in2_data = cst_2__icmp_9__data__0__anchor__in;
	assign cst_2__icmp_9__data__0__anchor__out = cst_2_out1_data;
	assign icmp_9_in2_valid = cst_2__icmp_9__valid__0__anchor__in;
	assign cst_2__icmp_9__valid__0__anchor__out = cst_2_out1_valid;
	assign cst_2_out1_ready = cst_2__icmp_9__ready__0__anchor__in;
	assign cst_2__icmp_9__ready__0__anchor__out = icmp_9_in2_ready;
	assign icmp_9_clk = clk;
	assign icmp_9_rst = rst;
	assign fork_16_in1_data = icmp_9__fork_16__data__0__anchor__in;
	assign icmp_9__fork_16__data__0__anchor__out = icmp_9_out1_data;
	assign fork_16_in1_valid = icmp_9__fork_16__valid__0__anchor__in;
	assign icmp_9__fork_16__valid__0__anchor__out = icmp_9_out1_valid;
	assign icmp_9_out1_ready = icmp_9__fork_16__ready__0__anchor__in;
	assign icmp_9__fork_16__ready__0__anchor__out = fork_16_in1_ready;
	assign cst_3_clk = clk;
	assign cst_3_rst = rst;
	assign add_11_in2_data = cst_3__add_11__data__0__anchor__in;
	assign cst_3__add_11__data__0__anchor__out = cst_3_out1_data;
	assign add_11_in2_valid = cst_3__add_11__valid__0__anchor__in;
	assign cst_3__add_11__valid__0__anchor__out = cst_3_out1_valid;
	assign cst_3_out1_ready = cst_3__add_11__ready__0__anchor__in;
	assign cst_3__add_11__ready__0__anchor__out = add_11_in2_ready;
	assign add_11_clk = clk;
	assign add_11_rst = rst;
	assign load_14_in2_data = add_11__load_14__data__0__anchor__in;
	assign add_11__load_14__data__0__anchor__out = add_11_out1_data;
	assign load_14_in2_valid = add_11__load_14__valid__0__anchor__in;
	assign add_11__load_14__valid__0__anchor__out = add_11_out1_valid;
	assign add_11_out1_ready = add_11__load_14__ready__0__anchor__in;
	assign add_11__load_14__ready__0__anchor__out = load_14_in2_ready;
	assign load_14_clk = clk;
	assign load_14_rst = rst;
	assign icmp_15_in1_data = load_14__icmp_15__data__0__anchor__in;
	assign load_14__icmp_15__data__0__anchor__out = load_14_out1_data;
	assign icmp_15_in1_valid = load_14__icmp_15__valid__0__anchor__in;
	assign load_14__icmp_15__valid__0__anchor__out = load_14_out1_valid;
	assign load_14_out1_ready = load_14__icmp_15__ready__0__anchor__in;
	assign load_14__icmp_15__ready__0__anchor__out = icmp_15_in1_ready;
	assign MC_A_in4_data = load_14__MC_A__data__0__anchor__in;
	assign load_14__MC_A__data__0__anchor__out = load_14_out2_data;
	assign MC_A_in4_valid = load_14__MC_A__valid__0__anchor__in;
	assign load_14__MC_A__valid__0__anchor__out = load_14_out2_valid;
	assign load_14_out2_ready = load_14__MC_A__ready__0__anchor__in;
	assign load_14__MC_A__ready__0__anchor__out = MC_A_in4_ready;
	assign icmp_15_clk = clk;
	assign icmp_15_rst = rst;
	assign Buffer_58_in1_data = icmp_15__Buffer_58__data__0__anchor__in;
	assign icmp_15__Buffer_58__data__0__anchor__out = icmp_15_out1_data;
	assign Buffer_58_in1_valid = icmp_15__Buffer_58__valid__0__anchor__in;
	assign icmp_15__Buffer_58__valid__0__anchor__out = icmp_15_out1_valid;
	assign icmp_15_out1_ready = icmp_15__Buffer_58__ready__0__anchor__in;
	assign icmp_15__Buffer_58__ready__0__anchor__out = Buffer_58_in1_ready;
	assign cst_4_clk = clk;
	assign cst_4_rst = rst;
	assign add_17_in2_data = cst_4__add_17__data__0__anchor__in;
	assign cst_4__add_17__data__0__anchor__out = cst_4_out1_data;
	assign add_17_in2_valid = cst_4__add_17__valid__0__anchor__in;
	assign cst_4__add_17__valid__0__anchor__out = cst_4_out1_valid;
	assign cst_4_out1_ready = cst_4__add_17__ready__0__anchor__in;
	assign cst_4__add_17__ready__0__anchor__out = add_17_in2_ready;
	assign add_17_clk = clk;
	assign add_17_rst = rst;
	assign load_20_in2_data = add_17__load_20__data__0__anchor__in;
	assign add_17__load_20__data__0__anchor__out = add_17_out1_data;
	assign load_20_in2_valid = add_17__load_20__valid__0__anchor__in;
	assign add_17__load_20__valid__0__anchor__out = add_17_out1_valid;
	assign add_17_out1_ready = add_17__load_20__ready__0__anchor__in;
	assign add_17__load_20__ready__0__anchor__out = load_20_in2_ready;
	assign load_20_clk = clk;
	assign load_20_rst = rst;
	assign store_0_in1_data = load_20__store_0__data__0__anchor__in;
	assign load_20__store_0__data__0__anchor__out = load_20_out1_data;
	assign store_0_in1_valid = load_20__store_0__valid__0__anchor__in;
	assign load_20__store_0__valid__0__anchor__out = load_20_out1_valid;
	assign load_20_out1_ready = load_20__store_0__ready__0__anchor__in;
	assign load_20__store_0__ready__0__anchor__out = store_0_in1_ready;
	assign MC_A_in5_data = load_20__MC_A__data__0__anchor__in;
	assign load_20__MC_A__data__0__anchor__out = load_20_out2_data;
	assign MC_A_in5_valid = load_20__MC_A__valid__0__anchor__in;
	assign load_20__MC_A__valid__0__anchor__out = load_20_out2_valid;
	assign load_20_out2_ready = load_20__MC_A__ready__0__anchor__in;
	assign load_20__MC_A__ready__0__anchor__out = MC_A_in5_ready;
	assign store_0_clk = clk;
	assign store_0_rst = rst;
	assign MC_A_in7_data = store_0__MC_A__data__0__anchor__in;
	assign store_0__MC_A__data__0__anchor__out = store_0_out1_data;
	assign MC_A_in7_valid = store_0__MC_A__valid__0__anchor__in;
	assign store_0__MC_A__valid__0__anchor__out = store_0_out1_valid;
	assign store_0_out1_ready = store_0__MC_A__ready__0__anchor__in;
	assign store_0__MC_A__ready__0__anchor__out = MC_A_in7_ready;
	assign MC_A_in6_data = store_0__MC_A__data__1__anchor__in;
	assign store_0__MC_A__data__1__anchor__out = store_0_out2_data;
	assign MC_A_in6_valid = store_0__MC_A__valid__1__anchor__in;
	assign store_0__MC_A__valid__1__anchor__out = store_0_out2_valid;
	assign store_0_out2_ready = store_0__MC_A__ready__1__anchor__in;
	assign store_0__MC_A__ready__1__anchor__out = MC_A_in6_ready;
	assign cst_5_clk = clk;
	assign cst_5_rst = rst;
	assign add_23_in2_data = cst_5__add_23__data__0__anchor__in;
	assign cst_5__add_23__data__0__anchor__out = cst_5_out1_data;
	assign add_23_in2_valid = cst_5__add_23__valid__0__anchor__in;
	assign cst_5__add_23__valid__0__anchor__out = cst_5_out1_valid;
	assign cst_5_out1_ready = cst_5__add_23__ready__0__anchor__in;
	assign cst_5__add_23__ready__0__anchor__out = add_23_in2_ready;
	assign add_23_clk = clk;
	assign add_23_rst = rst;
	assign branch_15_in1_data = add_23__branch_15__data__0__anchor__in;
	assign add_23__branch_15__data__0__anchor__out = add_23_out1_data;
	assign branch_15_in1_valid = add_23__branch_15__valid__0__anchor__in;
	assign add_23__branch_15__valid__0__anchor__out = add_23_out1_valid;
	assign add_23_out1_ready = add_23__branch_15__ready__0__anchor__in;
	assign add_23__branch_15__ready__0__anchor__out = branch_15_in1_ready;
	assign brCst_block6_clk = clk;
	assign brCst_block6_rst = rst;
	assign fork_18_in1_data = brCst_block6__fork_18__data__0__anchor__in;
	assign brCst_block6__fork_18__data__0__anchor__out = brCst_block6_out1_data;
	assign fork_18_in1_valid = brCst_block6__fork_18__valid__0__anchor__in;
	assign brCst_block6__fork_18__valid__0__anchor__out = brCst_block6_out1_valid;
	assign brCst_block6_out1_ready = brCst_block6__fork_18__ready__0__anchor__in;
	assign brCst_block6__fork_18__ready__0__anchor__out = fork_18_in1_ready;
	assign store_1_clk = clk;
	assign store_1_rst = rst;
	assign MC_A_in9_data = store_1__MC_A__data__0__anchor__in;
	assign store_1__MC_A__data__0__anchor__out = store_1_out1_data;
	assign MC_A_in9_valid = store_1__MC_A__valid__0__anchor__in;
	assign store_1__MC_A__valid__0__anchor__out = store_1_out1_valid;
	assign store_1_out1_ready = store_1__MC_A__ready__0__anchor__in;
	assign store_1__MC_A__ready__0__anchor__out = MC_A_in9_ready;
	assign MC_A_in8_data = store_1__MC_A__data__1__anchor__in;
	assign store_1__MC_A__data__1__anchor__out = store_1_out2_data;
	assign MC_A_in8_valid = store_1__MC_A__valid__1__anchor__in;
	assign store_1__MC_A__valid__1__anchor__out = store_1_out2_valid;
	assign store_1_out2_ready = store_1__MC_A__ready__1__anchor__in;
	assign store_1__MC_A__ready__1__anchor__out = MC_A_in8_ready;
	assign cst_6_clk = clk;
	assign cst_6_rst = rst;
	assign add_27_in2_data = cst_6__add_27__data__0__anchor__in;
	assign cst_6__add_27__data__0__anchor__out = cst_6_out1_data;
	assign add_27_in2_valid = cst_6__add_27__valid__0__anchor__in;
	assign cst_6__add_27__valid__0__anchor__out = cst_6_out1_valid;
	assign cst_6_out1_ready = cst_6__add_27__ready__0__anchor__in;
	assign cst_6__add_27__ready__0__anchor__out = add_27_in2_ready;
	assign add_27_clk = clk;
	assign add_27_rst = rst;
	assign fork_3_in1_data = add_27__fork_3__data__0__anchor__in;
	assign add_27__fork_3__data__0__anchor__out = add_27_out1_data;
	assign fork_3_in1_valid = add_27__fork_3__valid__0__anchor__in;
	assign add_27__fork_3__valid__0__anchor__out = add_27_out1_valid;
	assign add_27_out1_ready = add_27__fork_3__ready__0__anchor__in;
	assign add_27__fork_3__ready__0__anchor__out = fork_3_in1_ready;
	assign icmp_28_clk = clk;
	assign icmp_28_rst = rst;
	assign fork_19_in1_data = icmp_28__fork_19__data__0__anchor__in;
	assign icmp_28__fork_19__data__0__anchor__out = icmp_28_out1_data;
	assign fork_19_in1_valid = icmp_28__fork_19__valid__0__anchor__in;
	assign icmp_28__fork_19__valid__0__anchor__out = icmp_28_out1_valid;
	assign icmp_28_out1_ready = icmp_28__fork_19__ready__0__anchor__in;
	assign icmp_28__fork_19__ready__0__anchor__out = fork_19_in1_ready;
	assign ret_0_clk = clk;
	assign ret_0_rst = rst;
	assign end_0_in2_data = ret_0__end_0__data__0__anchor__in;
	assign ret_0__end_0__data__0__anchor__out = ret_0_out1_data;
	assign end_0_in2_valid = ret_0__end_0__valid__0__anchor__in;
	assign ret_0__end_0__valid__0__anchor__out = ret_0_out1_valid;
	assign ret_0_out1_ready = ret_0__end_0__ready__0__anchor__in;
	assign ret_0__end_0__ready__0__anchor__out = end_0_in2_ready;
	assign phi_n0_clk = clk;
	assign phi_n0_rst = rst;
	assign branch_2_in1_data = phi_n0__branch_2__data__0__anchor__in;
	assign phi_n0__branch_2__data__0__anchor__out = phi_n0_out1_data;
	assign branch_2_in1_valid = phi_n0__branch_2__valid__0__anchor__in;
	assign phi_n0__branch_2__valid__0__anchor__out = phi_n0_out1_valid;
	assign phi_n0_out1_ready = phi_n0__branch_2__ready__0__anchor__in;
	assign phi_n0__branch_2__ready__0__anchor__out = branch_2_in1_ready;
	assign phi_n1_clk = clk;
	assign phi_n1_rst = rst;
	assign branch_4_in1_data = phi_n1__branch_4__data__0__anchor__in;
	assign phi_n1__branch_4__data__0__anchor__out = phi_n1_out1_data;
	assign branch_4_in1_valid = phi_n1__branch_4__valid__0__anchor__in;
	assign phi_n1__branch_4__valid__0__anchor__out = phi_n1_out1_valid;
	assign phi_n1_out1_ready = phi_n1__branch_4__ready__0__anchor__in;
	assign phi_n1__branch_4__ready__0__anchor__out = branch_4_in1_ready;
	assign phi_n2_clk = clk;
	assign phi_n2_rst = rst;
	assign store_1_in1_data = phi_n2__store_1__data__0__anchor__in;
	assign phi_n2__store_1__data__0__anchor__out = phi_n2_out1_data;
	assign store_1_in1_valid = phi_n2__store_1__valid__0__anchor__in;
	assign phi_n2__store_1__valid__0__anchor__out = phi_n2_out1_valid;
	assign phi_n2_out1_ready = phi_n2__store_1__ready__0__anchor__in;
	assign phi_n2__store_1__ready__0__anchor__out = store_1_in1_ready;
	assign phi_n3_clk = clk;
	assign phi_n3_rst = rst;
	assign store_1_in2_data = phi_n3__store_1__data__0__anchor__in;
	assign phi_n3__store_1__data__0__anchor__out = phi_n3_out1_data;
	assign store_1_in2_valid = phi_n3__store_1__valid__0__anchor__in;
	assign phi_n3__store_1__valid__0__anchor__out = phi_n3_out1_valid;
	assign phi_n3_out1_ready = phi_n3__store_1__ready__0__anchor__in;
	assign phi_n3__store_1__ready__0__anchor__out = store_1_in2_ready;
	assign phi_n4_clk = clk;
	assign phi_n4_rst = rst;
	assign add_27_in1_data = phi_n4__add_27__data__0__anchor__in;
	assign phi_n4__add_27__data__0__anchor__out = phi_n4_out1_data;
	assign add_27_in1_valid = phi_n4__add_27__valid__0__anchor__in;
	assign phi_n4__add_27__valid__0__anchor__out = phi_n4_out1_valid;
	assign phi_n4_out1_ready = phi_n4__add_27__ready__0__anchor__in;
	assign phi_n4__add_27__ready__0__anchor__out = add_27_in1_ready;
	assign phi_n5_clk = clk;
	assign phi_n5_rst = rst;
	assign fork_4_in1_data = phi_n5__fork_4__data__0__anchor__in;
	assign phi_n5__fork_4__data__0__anchor__out = phi_n5_out1_data;
	assign fork_4_in1_valid = phi_n5__fork_4__valid__0__anchor__in;
	assign phi_n5__fork_4__valid__0__anchor__out = phi_n5_out1_valid;
	assign phi_n5_out1_ready = phi_n5__fork_4__ready__0__anchor__in;
	assign phi_n5__fork_4__ready__0__anchor__out = fork_4_in1_ready;
	assign phi_n6_clk = clk;
	assign phi_n6_rst = rst;
	assign branch_8_in1_data = phi_n6__branch_8__data__0__anchor__in;
	assign phi_n6__branch_8__data__0__anchor__out = phi_n6_out1_data;
	assign branch_8_in1_valid = phi_n6__branch_8__valid__0__anchor__in;
	assign phi_n6__branch_8__valid__0__anchor__out = phi_n6_out1_valid;
	assign phi_n6_out1_ready = phi_n6__branch_8__ready__0__anchor__in;
	assign phi_n6__branch_8__ready__0__anchor__out = branch_8_in1_ready;
	assign phi_n7_clk = clk;
	assign phi_n7_rst = rst;
	assign branch_9_in1_data = phi_n7__branch_9__data__0__anchor__in;
	assign phi_n7__branch_9__data__0__anchor__out = phi_n7_out1_data;
	assign branch_9_in1_valid = phi_n7__branch_9__valid__0__anchor__in;
	assign phi_n7__branch_9__valid__0__anchor__out = phi_n7_out1_valid;
	assign phi_n7_out1_ready = phi_n7__branch_9__ready__0__anchor__in;
	assign phi_n7__branch_9__ready__0__anchor__out = branch_9_in1_ready;
	assign phi_n8_clk = clk;
	assign phi_n8_rst = rst;
	assign branch_10_in1_data = phi_n8__branch_10__data__0__anchor__in;
	assign phi_n8__branch_10__data__0__anchor__out = phi_n8_out1_data;
	assign branch_10_in1_valid = phi_n8__branch_10__valid__0__anchor__in;
	assign phi_n8__branch_10__valid__0__anchor__out = phi_n8_out1_valid;
	assign phi_n8_out1_ready = phi_n8__branch_10__ready__0__anchor__in;
	assign phi_n8__branch_10__ready__0__anchor__out = branch_10_in1_ready;
	assign phi_n9_clk = clk;
	assign phi_n9_rst = rst;
	assign fork_8_in1_data = phi_n9__fork_8__data__0__anchor__in;
	assign phi_n9__fork_8__data__0__anchor__out = phi_n9_out1_data;
	assign fork_8_in1_valid = phi_n9__fork_8__valid__0__anchor__in;
	assign phi_n9__fork_8__valid__0__anchor__out = phi_n9_out1_valid;
	assign phi_n9_out1_ready = phi_n9__fork_8__ready__0__anchor__in;
	assign phi_n9__fork_8__ready__0__anchor__out = fork_8_in1_ready;
	assign phi_n10_clk = clk;
	assign phi_n10_rst = rst;
	assign branch_16_in1_data = phi_n10__branch_16__data__0__anchor__in;
	assign phi_n10__branch_16__data__0__anchor__out = phi_n10_out1_data;
	assign branch_16_in1_valid = phi_n10__branch_16__valid__0__anchor__in;
	assign phi_n10__branch_16__valid__0__anchor__out = phi_n10_out1_valid;
	assign phi_n10_out1_ready = phi_n10__branch_16__ready__0__anchor__in;
	assign phi_n10__branch_16__ready__0__anchor__out = branch_16_in1_ready;
	assign phi_n11_clk = clk;
	assign phi_n11_rst = rst;
	assign branch_17_in1_data = phi_n11__branch_17__data__0__anchor__in;
	assign phi_n11__branch_17__data__0__anchor__out = phi_n11_out1_data;
	assign branch_17_in1_valid = phi_n11__branch_17__valid__0__anchor__in;
	assign phi_n11__branch_17__valid__0__anchor__out = phi_n11_out1_valid;
	assign phi_n11_out1_ready = phi_n11__branch_17__ready__0__anchor__in;
	assign phi_n11__branch_17__ready__0__anchor__out = branch_17_in1_ready;
	assign phi_n12_clk = clk;
	assign phi_n12_rst = rst;
	assign branch_18_in1_data = phi_n12__branch_18__data__0__anchor__in;
	assign phi_n12__branch_18__data__0__anchor__out = phi_n12_out1_data;
	assign branch_18_in1_valid = phi_n12__branch_18__valid__0__anchor__in;
	assign phi_n12__branch_18__valid__0__anchor__out = phi_n12_out1_valid;
	assign phi_n12_out1_ready = phi_n12__branch_18__ready__0__anchor__in;
	assign phi_n12__branch_18__ready__0__anchor__out = branch_18_in1_ready;
	assign phi_n13_clk = clk;
	assign phi_n13_rst = rst;
	assign fork_9_in1_data = phi_n13__fork_9__data__0__anchor__in;
	assign phi_n13__fork_9__data__0__anchor__out = phi_n13_out1_data;
	assign fork_9_in1_valid = phi_n13__fork_9__valid__0__anchor__in;
	assign phi_n13__fork_9__valid__0__anchor__out = phi_n13_out1_valid;
	assign phi_n13_out1_ready = phi_n13__fork_9__ready__0__anchor__in;
	assign phi_n13__fork_9__ready__0__anchor__out = fork_9_in1_ready;
	assign phi_n14_clk = clk;
	assign phi_n14_rst = rst;
	assign fork_10_in1_data = phi_n14__fork_10__data__0__anchor__in;
	assign phi_n14__fork_10__data__0__anchor__out = phi_n14_out1_data;
	assign fork_10_in1_valid = phi_n14__fork_10__valid__0__anchor__in;
	assign phi_n14__fork_10__valid__0__anchor__out = phi_n14_out1_valid;
	assign phi_n14_out1_ready = phi_n14__fork_10__ready__0__anchor__in;
	assign phi_n14__fork_10__ready__0__anchor__out = fork_10_in1_ready;
	assign phi_n15_clk = clk;
	assign phi_n15_rst = rst;
	assign branch_13_in1_data = phi_n15__branch_13__data__0__anchor__in;
	assign phi_n15__branch_13__data__0__anchor__out = phi_n15_out1_data;
	assign branch_13_in1_valid = phi_n15__branch_13__valid__0__anchor__in;
	assign phi_n15__branch_13__valid__0__anchor__out = phi_n15_out1_valid;
	assign phi_n15_out1_ready = phi_n15__branch_13__ready__0__anchor__in;
	assign phi_n15__branch_13__ready__0__anchor__out = branch_13_in1_ready;
	assign phi_n16_clk = clk;
	assign phi_n16_rst = rst;
	assign branch_14_in1_data = phi_n16__branch_14__data__0__anchor__in;
	assign phi_n16__branch_14__data__0__anchor__out = phi_n16_out1_data;
	assign branch_14_in1_valid = phi_n16__branch_14__valid__0__anchor__in;
	assign phi_n16__branch_14__valid__0__anchor__out = phi_n16_out1_valid;
	assign phi_n16_out1_ready = phi_n16__branch_14__ready__0__anchor__in;
	assign phi_n16__branch_14__ready__0__anchor__out = branch_14_in1_ready;
	assign fork_0_clk = clk;
	assign fork_0_rst = rst;
	assign icmp_0_in1_data = fork_0__icmp_0__data__0__anchor__in;
	assign fork_0__icmp_0__data__0__anchor__out = fork_0_out1_data;
	assign icmp_0_in1_valid = fork_0__icmp_0__valid__0__anchor__in;
	assign fork_0__icmp_0__valid__0__anchor__out = fork_0_out1_valid;
	assign fork_0_out1_ready = fork_0__icmp_0__ready__0__anchor__in;
	assign fork_0__icmp_0__ready__0__anchor__out = icmp_0_in1_ready;
	assign branch_0_in1_data = fork_0__branch_0__data__0__anchor__in;
	assign fork_0__branch_0__data__0__anchor__out = fork_0_out2_data;
	assign branch_0_in1_valid = fork_0__branch_0__valid__0__anchor__in;
	assign fork_0__branch_0__valid__0__anchor__out = fork_0_out2_valid;
	assign fork_0_out2_ready = fork_0__branch_0__ready__0__anchor__in;
	assign fork_0__branch_0__ready__0__anchor__out = branch_0_in1_ready;
	assign fork_1_clk = clk;
	assign fork_1_rst = rst;
	assign load_6_in2_data = fork_1__load_6__data__0__anchor__in;
	assign fork_1__load_6__data__0__anchor__out = fork_1_out1_data;
	assign load_6_in2_valid = fork_1__load_6__valid__0__anchor__in;
	assign fork_1__load_6__valid__0__anchor__out = fork_1_out1_valid;
	assign fork_1_out1_ready = fork_1__load_6__ready__0__anchor__in;
	assign fork_1__load_6__ready__0__anchor__out = load_6_in2_ready;
	assign branch_5_in1_data = fork_1__branch_5__data__0__anchor__in;
	assign fork_1__branch_5__data__0__anchor__out = fork_1_out2_data;
	assign branch_5_in1_valid = fork_1__branch_5__valid__0__anchor__in;
	assign fork_1__branch_5__valid__0__anchor__out = fork_1_out2_valid;
	assign fork_1_out2_ready = fork_1__branch_5__ready__0__anchor__in;
	assign fork_1__branch_5__ready__0__anchor__out = branch_5_in1_ready;
	assign branch_6_in1_data = fork_1__branch_6__data__0__anchor__in;
	assign fork_1__branch_6__data__0__anchor__out = fork_1_out3_data;
	assign branch_6_in1_valid = fork_1__branch_6__valid__0__anchor__in;
	assign fork_1__branch_6__valid__0__anchor__out = fork_1_out3_valid;
	assign fork_1_out3_ready = fork_1__branch_6__ready__0__anchor__in;
	assign fork_1__branch_6__ready__0__anchor__out = branch_6_in1_ready;
	assign fork_2_clk = clk;
	assign fork_2_rst = rst;
	assign icmp_9_in1_data = fork_2__icmp_9__data__0__anchor__in;
	assign fork_2__icmp_9__data__0__anchor__out = fork_2_out1_data;
	assign icmp_9_in1_valid = fork_2__icmp_9__valid__0__anchor__in;
	assign fork_2__icmp_9__valid__0__anchor__out = fork_2_out1_valid;
	assign fork_2_out1_ready = fork_2__icmp_9__ready__0__anchor__in;
	assign fork_2__icmp_9__ready__0__anchor__out = icmp_9_in1_ready;
	assign branch_7_in1_data = fork_2__branch_7__data__0__anchor__in;
	assign fork_2__branch_7__data__0__anchor__out = fork_2_out2_data;
	assign branch_7_in1_valid = fork_2__branch_7__valid__0__anchor__in;
	assign fork_2__branch_7__valid__0__anchor__out = fork_2_out2_valid;
	assign fork_2_out2_ready = fork_2__branch_7__ready__0__anchor__in;
	assign fork_2__branch_7__ready__0__anchor__out = branch_7_in1_ready;
	assign fork_3_clk = clk;
	assign fork_3_rst = rst;
	assign icmp_28_in1_data = fork_3__icmp_28__data__0__anchor__in;
	assign fork_3__icmp_28__data__0__anchor__out = fork_3_out1_data;
	assign icmp_28_in1_valid = fork_3__icmp_28__valid__0__anchor__in;
	assign fork_3__icmp_28__valid__0__anchor__out = fork_3_out1_valid;
	assign fork_3_out1_ready = fork_3__icmp_28__ready__0__anchor__in;
	assign fork_3__icmp_28__ready__0__anchor__out = icmp_28_in1_ready;
	assign branch_19_in1_data = fork_3__branch_19__data__0__anchor__in;
	assign fork_3__branch_19__data__0__anchor__out = fork_3_out2_data;
	assign branch_19_in1_valid = fork_3__branch_19__valid__0__anchor__in;
	assign fork_3__branch_19__valid__0__anchor__out = fork_3_out2_valid;
	assign fork_3_out2_ready = fork_3__branch_19__ready__0__anchor__in;
	assign fork_3__branch_19__ready__0__anchor__out = branch_19_in1_ready;
	assign fork_4_clk = clk;
	assign fork_4_rst = rst;
	assign icmp_28_in2_data = fork_4__icmp_28__data__0__anchor__in;
	assign fork_4__icmp_28__data__0__anchor__out = fork_4_out1_data;
	assign icmp_28_in2_valid = fork_4__icmp_28__valid__0__anchor__in;
	assign fork_4__icmp_28__valid__0__anchor__out = fork_4_out1_valid;
	assign fork_4_out1_ready = fork_4__icmp_28__ready__0__anchor__in;
	assign fork_4__icmp_28__ready__0__anchor__out = icmp_28_in2_ready;
	assign branch_20_in1_data = fork_4__branch_20__data__0__anchor__in;
	assign fork_4__branch_20__data__0__anchor__out = fork_4_out2_data;
	assign branch_20_in1_valid = fork_4__branch_20__valid__0__anchor__in;
	assign fork_4__branch_20__valid__0__anchor__out = fork_4_out2_valid;
	assign fork_4_out2_ready = fork_4__branch_20__ready__0__anchor__in;
	assign fork_4__branch_20__ready__0__anchor__out = branch_20_in1_ready;
	assign fork_8_clk = clk;
	assign fork_8_rst = rst;
	assign add_17_in1_data = fork_8__add_17__data__0__anchor__in;
	assign fork_8__add_17__data__0__anchor__out = fork_8_out1_data;
	assign add_17_in1_valid = fork_8__add_17__valid__0__anchor__in;
	assign fork_8__add_17__valid__0__anchor__out = fork_8_out1_valid;
	assign fork_8_out1_ready = fork_8__add_17__ready__0__anchor__in;
	assign fork_8__add_17__ready__0__anchor__out = add_17_in1_ready;
	assign store_0_in2_data = fork_8__store_0__data__0__anchor__in;
	assign fork_8__store_0__data__0__anchor__out = fork_8_out2_data;
	assign store_0_in2_valid = fork_8__store_0__valid__0__anchor__in;
	assign fork_8__store_0__valid__0__anchor__out = fork_8_out2_valid;
	assign fork_8_out2_ready = fork_8__store_0__ready__0__anchor__in;
	assign fork_8__store_0__ready__0__anchor__out = store_0_in2_ready;
	assign add_23_in1_data = fork_8__add_23__data__0__anchor__in;
	assign fork_8__add_23__data__0__anchor__out = fork_8_out3_data;
	assign add_23_in1_valid = fork_8__add_23__valid__0__anchor__in;
	assign fork_8__add_23__valid__0__anchor__out = fork_8_out3_valid;
	assign fork_8_out3_ready = fork_8__add_23__ready__0__anchor__in;
	assign fork_8__add_23__ready__0__anchor__out = add_23_in1_ready;
	assign fork_9_clk = clk;
	assign fork_9_rst = rst;
	assign add_11_in1_data = fork_9__add_11__data__0__anchor__in;
	assign fork_9__add_11__data__0__anchor__out = fork_9_out1_data;
	assign add_11_in1_valid = fork_9__add_11__valid__0__anchor__in;
	assign fork_9__add_11__valid__0__anchor__out = fork_9_out1_valid;
	assign fork_9_out1_ready = fork_9__add_11__ready__0__anchor__in;
	assign fork_9__add_11__ready__0__anchor__out = add_11_in1_ready;
	assign branch_11_in1_data = fork_9__branch_11__data__0__anchor__in;
	assign fork_9__branch_11__data__0__anchor__out = fork_9_out2_data;
	assign branch_11_in1_valid = fork_9__branch_11__valid__0__anchor__in;
	assign fork_9__branch_11__valid__0__anchor__out = fork_9_out2_valid;
	assign fork_9_out2_ready = fork_9__branch_11__ready__0__anchor__in;
	assign fork_9__branch_11__ready__0__anchor__out = branch_11_in1_ready;
	assign fork_10_clk = clk;
	assign fork_10_rst = rst;
	assign icmp_15_in2_data = fork_10__icmp_15__data__0__anchor__in;
	assign fork_10__icmp_15__data__0__anchor__out = fork_10_out1_data;
	assign icmp_15_in2_valid = fork_10__icmp_15__valid__0__anchor__in;
	assign fork_10__icmp_15__valid__0__anchor__out = fork_10_out1_valid;
	assign fork_10_out1_ready = fork_10__icmp_15__ready__0__anchor__in;
	assign fork_10__icmp_15__ready__0__anchor__out = icmp_15_in2_ready;
	assign branch_12_in1_data = fork_10__branch_12__data__0__anchor__in;
	assign fork_10__branch_12__data__0__anchor__out = fork_10_out2_data;
	assign branch_12_in1_valid = fork_10__branch_12__valid__0__anchor__in;
	assign fork_10__branch_12__valid__0__anchor__out = fork_10_out2_valid;
	assign fork_10_out2_ready = fork_10__branch_12__ready__0__anchor__in;
	assign fork_10__branch_12__ready__0__anchor__out = branch_12_in1_ready;
	assign branch_0_clk = clk;
	assign branch_0_rst = rst;
	assign sink_0_in1_data = branch_0__sink_0__data__0__anchor__in;
	assign branch_0__sink_0__data__0__anchor__out = branch_0_out1_data;
	assign sink_0_in1_valid = branch_0__sink_0__valid__0__anchor__in;
	assign branch_0__sink_0__valid__0__anchor__out = branch_0_out1_valid;
	assign branch_0_out1_ready = branch_0__sink_0__ready__0__anchor__in;
	assign branch_0__sink_0__ready__0__anchor__out = sink_0_in1_ready;
	assign phi_n0_in1_data = branch_0__phi_n0__data__0__anchor__in;
	assign branch_0__phi_n0__data__0__anchor__out = branch_0_out2_data;
	assign phi_n0_in1_valid = branch_0__phi_n0__valid__0__anchor__in;
	assign branch_0__phi_n0__valid__0__anchor__out = branch_0_out2_valid;
	assign branch_0_out2_ready = branch_0__phi_n0__ready__0__anchor__in;
	assign branch_0__phi_n0__ready__0__anchor__out = phi_n0_in1_ready;
	assign branch_1_clk = clk;
	assign branch_1_rst = rst;
	assign phi_3_in2_data = branch_1__phi_3__data__0__anchor__in;
	assign branch_1__phi_3__data__0__anchor__out = branch_1_out1_data;
	assign phi_3_in2_valid = branch_1__phi_3__valid__0__anchor__in;
	assign branch_1__phi_3__valid__0__anchor__out = branch_1_out1_valid;
	assign branch_1_out1_ready = branch_1__phi_3__ready__0__anchor__in;
	assign branch_1__phi_3__ready__0__anchor__out = phi_3_in2_ready;
	assign sink_1_in1_data = branch_1__sink_1__data__0__anchor__in;
	assign branch_1__sink_1__data__0__anchor__out = branch_1_out2_data;
	assign sink_1_in1_valid = branch_1__sink_1__valid__0__anchor__in;
	assign branch_1__sink_1__valid__0__anchor__out = branch_1_out2_valid;
	assign branch_1_out2_ready = branch_1__sink_1__ready__0__anchor__in;
	assign branch_1__sink_1__ready__0__anchor__out = sink_1_in1_ready;
	assign branch_2_clk = clk;
	assign branch_2_rst = rst;
	assign phi_n1_in1_data = branch_2__phi_n1__data__0__anchor__in;
	assign branch_2__phi_n1__data__0__anchor__out = branch_2_out1_data;
	assign phi_n1_in1_valid = branch_2__phi_n1__valid__0__anchor__in;
	assign branch_2__phi_n1__valid__0__anchor__out = branch_2_out1_valid;
	assign branch_2_out1_ready = branch_2__phi_n1__ready__0__anchor__in;
	assign branch_2__phi_n1__ready__0__anchor__out = phi_n1_in1_ready;
	assign sink_2_in1_data = branch_2__sink_2__data__0__anchor__in;
	assign branch_2__sink_2__data__0__anchor__out = branch_2_out2_data;
	assign sink_2_in1_valid = branch_2__sink_2__valid__0__anchor__in;
	assign branch_2__sink_2__valid__0__anchor__out = branch_2_out2_valid;
	assign branch_2_out2_ready = branch_2__sink_2__ready__0__anchor__in;
	assign branch_2__sink_2__ready__0__anchor__out = sink_2_in1_ready;
	assign fork_14_clk = clk;
	assign fork_14_rst = rst;
	assign branch_2_in2_data = fork_14__branch_2__data__0__anchor__in;
	assign fork_14__branch_2__data__0__anchor__out = fork_14_out1_data;
	assign branch_2_in2_valid = fork_14__branch_2__valid__0__anchor__in;
	assign fork_14__branch_2__valid__0__anchor__out = fork_14_out1_valid;
	assign fork_14_out1_ready = fork_14__branch_2__ready__0__anchor__in;
	assign fork_14__branch_2__ready__0__anchor__out = branch_2_in2_ready;
	assign branch_1_in2_data = fork_14__branch_1__data__0__anchor__in;
	assign fork_14__branch_1__data__0__anchor__out = fork_14_out2_data;
	assign branch_1_in2_valid = fork_14__branch_1__valid__0__anchor__in;
	assign fork_14__branch_1__valid__0__anchor__out = fork_14_out2_valid;
	assign fork_14_out2_ready = fork_14__branch_1__ready__0__anchor__in;
	assign fork_14__branch_1__ready__0__anchor__out = branch_1_in2_ready;
	assign branchC_22_in2_data = fork_14__branchC_22__data__0__anchor__in;
	assign fork_14__branchC_22__data__0__anchor__out = fork_14_out3_data;
	assign branchC_22_in2_valid = fork_14__branchC_22__valid__0__anchor__in;
	assign fork_14__branchC_22__valid__0__anchor__out = fork_14_out3_valid;
	assign fork_14_out3_ready = fork_14__branchC_22__ready__0__anchor__in;
	assign fork_14__branchC_22__ready__0__anchor__out = branchC_22_in2_ready;
	assign branch_3_clk = clk;
	assign branch_3_rst = rst;
	assign phi_n6_in1_data = branch_3__phi_n6__data__0__anchor__in;
	assign branch_3__phi_n6__data__0__anchor__out = branch_3_out1_data;
	assign phi_n6_in1_valid = branch_3__phi_n6__valid__0__anchor__in;
	assign branch_3__phi_n6__valid__0__anchor__out = branch_3_out1_valid;
	assign branch_3_out1_ready = branch_3__phi_n6__ready__0__anchor__in;
	assign branch_3__phi_n6__ready__0__anchor__out = phi_n6_in1_ready;
	assign sink_3_in1_data = branch_3__sink_3__data__0__anchor__in;
	assign branch_3__sink_3__data__0__anchor__out = branch_3_out2_data;
	assign sink_3_in1_valid = branch_3__sink_3__valid__0__anchor__in;
	assign branch_3__sink_3__valid__0__anchor__out = branch_3_out2_valid;
	assign branch_3_out2_ready = branch_3__sink_3__ready__0__anchor__in;
	assign branch_3__sink_3__ready__0__anchor__out = sink_3_in1_ready;
	assign branch_4_clk = clk;
	assign branch_4_rst = rst;
	assign phi_n8_in1_data = branch_4__phi_n8__data__0__anchor__in;
	assign branch_4__phi_n8__data__0__anchor__out = branch_4_out1_data;
	assign phi_n8_in1_valid = branch_4__phi_n8__valid__0__anchor__in;
	assign branch_4__phi_n8__valid__0__anchor__out = branch_4_out1_valid;
	assign branch_4_out1_ready = branch_4__phi_n8__ready__0__anchor__in;
	assign branch_4__phi_n8__ready__0__anchor__out = phi_n8_in1_ready;
	assign sink_4_in1_data = branch_4__sink_4__data__0__anchor__in;
	assign branch_4__sink_4__data__0__anchor__out = branch_4_out2_data;
	assign sink_4_in1_valid = branch_4__sink_4__valid__0__anchor__in;
	assign branch_4__sink_4__valid__0__anchor__out = branch_4_out2_valid;
	assign branch_4_out2_ready = branch_4__sink_4__ready__0__anchor__in;
	assign branch_4__sink_4__ready__0__anchor__out = sink_4_in1_ready;
	assign branch_5_clk = clk;
	assign branch_5_rst = rst;
	assign phi_n7_in1_data = branch_5__phi_n7__data__0__anchor__in;
	assign branch_5__phi_n7__data__0__anchor__out = branch_5_out1_data;
	assign phi_n7_in1_valid = branch_5__phi_n7__valid__0__anchor__in;
	assign branch_5__phi_n7__valid__0__anchor__out = branch_5_out1_valid;
	assign branch_5_out1_ready = branch_5__phi_n7__ready__0__anchor__in;
	assign branch_5__phi_n7__ready__0__anchor__out = phi_n7_in1_ready;
	assign sink_5_in1_data = branch_5__sink_5__data__0__anchor__in;
	assign branch_5__sink_5__data__0__anchor__out = branch_5_out2_data;
	assign sink_5_in1_valid = branch_5__sink_5__valid__0__anchor__in;
	assign branch_5__sink_5__valid__0__anchor__out = branch_5_out2_valid;
	assign branch_5_out2_ready = branch_5__sink_5__ready__0__anchor__in;
	assign branch_5__sink_5__ready__0__anchor__out = sink_5_in1_ready;
	assign branch_6_clk = clk;
	assign branch_6_rst = rst;
	assign phi_8_in2_data = branch_6__phi_8__data__0__anchor__in;
	assign branch_6__phi_8__data__0__anchor__out = branch_6_out1_data;
	assign phi_8_in2_valid = branch_6__phi_8__valid__0__anchor__in;
	assign branch_6__phi_8__valid__0__anchor__out = branch_6_out1_valid;
	assign branch_6_out1_ready = branch_6__phi_8__ready__0__anchor__in;
	assign branch_6__phi_8__ready__0__anchor__out = phi_8_in2_ready;
	assign sink_6_in1_data = branch_6__sink_6__data__0__anchor__in;
	assign branch_6__sink_6__data__0__anchor__out = branch_6_out2_data;
	assign sink_6_in1_valid = branch_6__sink_6__valid__0__anchor__in;
	assign branch_6__sink_6__valid__0__anchor__out = branch_6_out2_valid;
	assign branch_6_out2_ready = branch_6__sink_6__ready__0__anchor__in;
	assign branch_6__sink_6__ready__0__anchor__out = sink_6_in1_ready;
	assign fork_15_clk = clk;
	assign fork_15_rst = rst;
	assign branch_6_in2_data = fork_15__branch_6__data__0__anchor__in;
	assign fork_15__branch_6__data__0__anchor__out = fork_15_out1_data;
	assign branch_6_in2_valid = fork_15__branch_6__valid__0__anchor__in;
	assign fork_15__branch_6__valid__0__anchor__out = fork_15_out1_valid;
	assign fork_15_out1_ready = fork_15__branch_6__ready__0__anchor__in;
	assign fork_15__branch_6__ready__0__anchor__out = branch_6_in2_ready;
	assign branch_5_in2_data = fork_15__branch_5__data__0__anchor__in;
	assign fork_15__branch_5__data__0__anchor__out = fork_15_out2_data;
	assign branch_5_in2_valid = fork_15__branch_5__valid__0__anchor__in;
	assign fork_15__branch_5__valid__0__anchor__out = fork_15_out2_valid;
	assign fork_15_out2_ready = fork_15__branch_5__ready__0__anchor__in;
	assign fork_15__branch_5__ready__0__anchor__out = branch_5_in2_ready;
	assign branch_4_in2_data = fork_15__branch_4__data__0__anchor__in;
	assign fork_15__branch_4__data__0__anchor__out = fork_15_out3_data;
	assign branch_4_in2_valid = fork_15__branch_4__valid__0__anchor__in;
	assign fork_15__branch_4__valid__0__anchor__out = fork_15_out3_valid;
	assign fork_15_out3_ready = fork_15__branch_4__ready__0__anchor__in;
	assign fork_15__branch_4__ready__0__anchor__out = branch_4_in2_ready;
	assign branch_3_in2_data = fork_15__branch_3__data__0__anchor__in;
	assign fork_15__branch_3__data__0__anchor__out = fork_15_out4_data;
	assign branch_3_in2_valid = fork_15__branch_3__valid__0__anchor__in;
	assign fork_15__branch_3__valid__0__anchor__out = fork_15_out4_valid;
	assign fork_15_out4_ready = fork_15__branch_3__ready__0__anchor__in;
	assign fork_15__branch_3__ready__0__anchor__out = branch_3_in2_ready;
	assign branchC_23_in2_data = fork_15__branchC_23__data__0__anchor__in;
	assign fork_15__branchC_23__data__0__anchor__out = fork_15_out5_data;
	assign branchC_23_in2_valid = fork_15__branchC_23__valid__0__anchor__in;
	assign fork_15__branchC_23__valid__0__anchor__out = fork_15_out5_valid;
	assign fork_15_out5_ready = fork_15__branchC_23__ready__0__anchor__in;
	assign fork_15__branchC_23__ready__0__anchor__out = branchC_23_in2_ready;
	assign branch_7_clk = clk;
	assign branch_7_rst = rst;
	assign phi_n13_in1_data = branch_7__phi_n13__data__0__anchor__in;
	assign branch_7__phi_n13__data__0__anchor__out = branch_7_out1_data;
	assign phi_n13_in1_valid = branch_7__phi_n13__valid__0__anchor__in;
	assign branch_7__phi_n13__valid__0__anchor__out = branch_7_out1_valid;
	assign branch_7_out1_ready = branch_7__phi_n13__ready__0__anchor__in;
	assign branch_7__phi_n13__ready__0__anchor__out = phi_n13_in1_ready;
	assign phi_n3_in1_data = branch_7__phi_n3__data__0__anchor__in;
	assign branch_7__phi_n3__data__0__anchor__out = branch_7_out2_data;
	assign phi_n3_in1_valid = branch_7__phi_n3__valid__0__anchor__in;
	assign branch_7__phi_n3__valid__0__anchor__out = branch_7_out2_valid;
	assign branch_7_out2_ready = branch_7__phi_n3__ready__0__anchor__in;
	assign branch_7__phi_n3__ready__0__anchor__out = phi_n3_in1_ready;
	assign branch_8_clk = clk;
	assign branch_8_rst = rst;
	assign phi_n14_in1_data = branch_8__phi_n14__data__0__anchor__in;
	assign branch_8__phi_n14__data__0__anchor__out = branch_8_out1_data;
	assign phi_n14_in1_valid = branch_8__phi_n14__valid__0__anchor__in;
	assign branch_8__phi_n14__valid__0__anchor__out = branch_8_out1_valid;
	assign branch_8_out1_ready = branch_8__phi_n14__ready__0__anchor__in;
	assign branch_8__phi_n14__ready__0__anchor__out = phi_n14_in1_ready;
	assign phi_n2_in1_data = branch_8__phi_n2__data__0__anchor__in;
	assign branch_8__phi_n2__data__0__anchor__out = branch_8_out2_data;
	assign phi_n2_in1_valid = branch_8__phi_n2__valid__0__anchor__in;
	assign branch_8__phi_n2__valid__0__anchor__out = branch_8_out2_valid;
	assign branch_8_out2_ready = branch_8__phi_n2__ready__0__anchor__in;
	assign branch_8__phi_n2__ready__0__anchor__out = phi_n2_in1_ready;
	assign branch_9_clk = clk;
	assign branch_9_rst = rst;
	assign phi_n15_in1_data = branch_9__phi_n15__data__0__anchor__in;
	assign branch_9__phi_n15__data__0__anchor__out = branch_9_out1_data;
	assign phi_n15_in1_valid = branch_9__phi_n15__valid__0__anchor__in;
	assign branch_9__phi_n15__valid__0__anchor__out = branch_9_out1_valid;
	assign branch_9_out1_ready = branch_9__phi_n15__ready__0__anchor__in;
	assign branch_9__phi_n15__ready__0__anchor__out = phi_n15_in1_ready;
	assign phi_n4_in1_data = branch_9__phi_n4__data__0__anchor__in;
	assign branch_9__phi_n4__data__0__anchor__out = branch_9_out2_data;
	assign phi_n4_in1_valid = branch_9__phi_n4__valid__0__anchor__in;
	assign branch_9__phi_n4__valid__0__anchor__out = branch_9_out2_valid;
	assign branch_9_out2_ready = branch_9__phi_n4__ready__0__anchor__in;
	assign branch_9__phi_n4__ready__0__anchor__out = phi_n4_in1_ready;
	assign branch_10_clk = clk;
	assign branch_10_rst = rst;
	assign phi_n16_in1_data = branch_10__phi_n16__data__0__anchor__in;
	assign branch_10__phi_n16__data__0__anchor__out = branch_10_out1_data;
	assign phi_n16_in1_valid = branch_10__phi_n16__valid__0__anchor__in;
	assign branch_10__phi_n16__valid__0__anchor__out = branch_10_out1_valid;
	assign branch_10_out1_ready = branch_10__phi_n16__ready__0__anchor__in;
	assign branch_10__phi_n16__ready__0__anchor__out = phi_n16_in1_ready;
	assign phi_n5_in1_data = branch_10__phi_n5__data__0__anchor__in;
	assign branch_10__phi_n5__data__0__anchor__out = branch_10_out2_data;
	assign phi_n5_in1_valid = branch_10__phi_n5__valid__0__anchor__in;
	assign branch_10__phi_n5__valid__0__anchor__out = branch_10_out2_valid;
	assign branch_10_out2_ready = branch_10__phi_n5__ready__0__anchor__in;
	assign branch_10__phi_n5__ready__0__anchor__out = phi_n5_in1_ready;
	assign fork_16_clk = clk;
	assign fork_16_rst = rst;
	assign branch_10_in2_data = fork_16__branch_10__data__0__anchor__in;
	assign fork_16__branch_10__data__0__anchor__out = fork_16_out1_data;
	assign branch_10_in2_valid = fork_16__branch_10__valid__0__anchor__in;
	assign fork_16__branch_10__valid__0__anchor__out = fork_16_out1_valid;
	assign fork_16_out1_ready = fork_16__branch_10__ready__0__anchor__in;
	assign fork_16__branch_10__ready__0__anchor__out = branch_10_in2_ready;
	assign branch_9_in2_data = fork_16__branch_9__data__0__anchor__in;
	assign fork_16__branch_9__data__0__anchor__out = fork_16_out2_data;
	assign branch_9_in2_valid = fork_16__branch_9__valid__0__anchor__in;
	assign fork_16__branch_9__valid__0__anchor__out = fork_16_out2_valid;
	assign fork_16_out2_ready = fork_16__branch_9__ready__0__anchor__in;
	assign fork_16__branch_9__ready__0__anchor__out = branch_9_in2_ready;
	assign branch_8_in2_data = fork_16__branch_8__data__0__anchor__in;
	assign fork_16__branch_8__data__0__anchor__out = fork_16_out3_data;
	assign branch_8_in2_valid = fork_16__branch_8__valid__0__anchor__in;
	assign fork_16__branch_8__valid__0__anchor__out = fork_16_out3_valid;
	assign fork_16_out3_ready = fork_16__branch_8__ready__0__anchor__in;
	assign fork_16__branch_8__ready__0__anchor__out = branch_8_in2_ready;
	assign branch_7_in2_data = fork_16__branch_7__data__0__anchor__in;
	assign fork_16__branch_7__data__0__anchor__out = fork_16_out4_data;
	assign branch_7_in2_valid = fork_16__branch_7__valid__0__anchor__in;
	assign fork_16__branch_7__valid__0__anchor__out = fork_16_out4_valid;
	assign fork_16_out4_ready = fork_16__branch_7__ready__0__anchor__in;
	assign fork_16__branch_7__ready__0__anchor__out = branch_7_in2_ready;
	assign branchC_24_in2_data = fork_16__branchC_24__data__0__anchor__in;
	assign fork_16__branchC_24__data__0__anchor__out = fork_16_out5_data;
	assign branchC_24_in2_valid = fork_16__branchC_24__valid__0__anchor__in;
	assign fork_16__branchC_24__valid__0__anchor__out = fork_16_out5_valid;
	assign fork_16_out5_ready = fork_16__branchC_24__ready__0__anchor__in;
	assign fork_16__branchC_24__ready__0__anchor__out = branchC_24_in2_ready;
	assign branch_11_clk = clk;
	assign branch_11_rst = rst;
	assign phi_n9_in1_data = branch_11__phi_n9__data__0__anchor__in;
	assign branch_11__phi_n9__data__0__anchor__out = branch_11_out1_data;
	assign phi_n9_in1_valid = branch_11__phi_n9__valid__0__anchor__in;
	assign branch_11__phi_n9__valid__0__anchor__out = branch_11_out1_valid;
	assign branch_11_out1_ready = branch_11__phi_n9__ready__0__anchor__in;
	assign branch_11__phi_n9__ready__0__anchor__out = phi_n9_in1_ready;
	assign phi_n3_in2_data = branch_11__phi_n3__data__0__anchor__in;
	assign branch_11__phi_n3__data__0__anchor__out = branch_11_out2_data;
	assign phi_n3_in2_valid = branch_11__phi_n3__valid__0__anchor__in;
	assign branch_11__phi_n3__valid__0__anchor__out = branch_11_out2_valid;
	assign branch_11_out2_ready = branch_11__phi_n3__ready__0__anchor__in;
	assign branch_11__phi_n3__ready__0__anchor__out = phi_n3_in2_ready;
	assign branch_12_clk = clk;
	assign branch_12_rst = rst;
	assign phi_n10_in1_data = branch_12__phi_n10__data__0__anchor__in;
	assign branch_12__phi_n10__data__0__anchor__out = branch_12_out1_data;
	assign phi_n10_in1_valid = branch_12__phi_n10__valid__0__anchor__in;
	assign branch_12__phi_n10__valid__0__anchor__out = branch_12_out1_valid;
	assign branch_12_out1_ready = branch_12__phi_n10__ready__0__anchor__in;
	assign branch_12__phi_n10__ready__0__anchor__out = phi_n10_in1_ready;
	assign phi_n2_in2_data = branch_12__phi_n2__data__0__anchor__in;
	assign branch_12__phi_n2__data__0__anchor__out = branch_12_out2_data;
	assign phi_n2_in2_valid = branch_12__phi_n2__valid__0__anchor__in;
	assign branch_12__phi_n2__valid__0__anchor__out = branch_12_out2_valid;
	assign branch_12_out2_ready = branch_12__phi_n2__ready__0__anchor__in;
	assign branch_12__phi_n2__ready__0__anchor__out = phi_n2_in2_ready;
	assign branch_13_clk = clk;
	assign branch_13_rst = rst;
	assign phi_n11_in1_data = branch_13__phi_n11__data__0__anchor__in;
	assign branch_13__phi_n11__data__0__anchor__out = branch_13_out1_data;
	assign phi_n11_in1_valid = branch_13__phi_n11__valid__0__anchor__in;
	assign branch_13__phi_n11__valid__0__anchor__out = branch_13_out1_valid;
	assign branch_13_out1_ready = branch_13__phi_n11__ready__0__anchor__in;
	assign branch_13__phi_n11__ready__0__anchor__out = phi_n11_in1_ready;
	assign phi_n4_in2_data = branch_13__phi_n4__data__0__anchor__in;
	assign branch_13__phi_n4__data__0__anchor__out = branch_13_out2_data;
	assign phi_n4_in2_valid = branch_13__phi_n4__valid__0__anchor__in;
	assign branch_13__phi_n4__valid__0__anchor__out = branch_13_out2_valid;
	assign branch_13_out2_ready = branch_13__phi_n4__ready__0__anchor__in;
	assign branch_13__phi_n4__ready__0__anchor__out = phi_n4_in2_ready;
	assign branch_14_clk = clk;
	assign branch_14_rst = rst;
	assign phi_n12_in1_data = branch_14__phi_n12__data__0__anchor__in;
	assign branch_14__phi_n12__data__0__anchor__out = branch_14_out1_data;
	assign phi_n12_in1_valid = branch_14__phi_n12__valid__0__anchor__in;
	assign branch_14__phi_n12__valid__0__anchor__out = branch_14_out1_valid;
	assign branch_14_out1_ready = branch_14__phi_n12__ready__0__anchor__in;
	assign branch_14__phi_n12__ready__0__anchor__out = phi_n12_in1_ready;
	assign phi_n5_in2_data = branch_14__phi_n5__data__0__anchor__in;
	assign branch_14__phi_n5__data__0__anchor__out = branch_14_out2_data;
	assign phi_n5_in2_valid = branch_14__phi_n5__valid__0__anchor__in;
	assign branch_14__phi_n5__valid__0__anchor__out = branch_14_out2_valid;
	assign branch_14_out2_ready = branch_14__phi_n5__ready__0__anchor__in;
	assign branch_14__phi_n5__ready__0__anchor__out = phi_n5_in2_ready;
	assign fork_17_clk = clk;
	assign fork_17_rst = rst;
	assign branch_14_in2_data = fork_17__branch_14__data__0__anchor__in;
	assign fork_17__branch_14__data__0__anchor__out = fork_17_out1_data;
	assign branch_14_in2_valid = fork_17__branch_14__valid__0__anchor__in;
	assign fork_17__branch_14__valid__0__anchor__out = fork_17_out1_valid;
	assign fork_17_out1_ready = fork_17__branch_14__ready__0__anchor__in;
	assign fork_17__branch_14__ready__0__anchor__out = branch_14_in2_ready;
	assign branch_13_in2_data = fork_17__branch_13__data__0__anchor__in;
	assign fork_17__branch_13__data__0__anchor__out = fork_17_out2_data;
	assign branch_13_in2_valid = fork_17__branch_13__valid__0__anchor__in;
	assign fork_17__branch_13__valid__0__anchor__out = fork_17_out2_valid;
	assign fork_17_out2_ready = fork_17__branch_13__ready__0__anchor__in;
	assign fork_17__branch_13__ready__0__anchor__out = branch_13_in2_ready;
	assign branch_12_in2_data = fork_17__branch_12__data__0__anchor__in;
	assign fork_17__branch_12__data__0__anchor__out = fork_17_out3_data;
	assign branch_12_in2_valid = fork_17__branch_12__valid__0__anchor__in;
	assign fork_17__branch_12__valid__0__anchor__out = fork_17_out3_valid;
	assign fork_17_out3_ready = fork_17__branch_12__ready__0__anchor__in;
	assign fork_17__branch_12__ready__0__anchor__out = branch_12_in2_ready;
	assign branch_11_in2_data = fork_17__branch_11__data__0__anchor__in;
	assign fork_17__branch_11__data__0__anchor__out = fork_17_out4_data;
	assign branch_11_in2_valid = fork_17__branch_11__valid__0__anchor__in;
	assign fork_17__branch_11__valid__0__anchor__out = fork_17_out4_valid;
	assign fork_17_out4_ready = fork_17__branch_11__ready__0__anchor__in;
	assign fork_17__branch_11__ready__0__anchor__out = branch_11_in2_ready;
	assign branchC_25_in2_data = fork_17__branchC_25__data__0__anchor__in;
	assign fork_17__branchC_25__data__0__anchor__out = fork_17_out5_data;
	assign branchC_25_in2_valid = fork_17__branchC_25__valid__0__anchor__in;
	assign fork_17__branchC_25__valid__0__anchor__out = fork_17_out5_valid;
	assign fork_17_out5_ready = fork_17__branchC_25__ready__0__anchor__in;
	assign fork_17__branchC_25__ready__0__anchor__out = branchC_25_in2_ready;
	assign branch_15_clk = clk;
	assign branch_15_rst = rst;
	assign Buffer_51_in1_data = branch_15__Buffer_51__data__0__anchor__in;
	assign branch_15__Buffer_51__data__0__anchor__out = branch_15_out1_data;
	assign Buffer_51_in1_valid = branch_15__Buffer_51__valid__0__anchor__in;
	assign branch_15__Buffer_51__valid__0__anchor__out = branch_15_out1_valid;
	assign branch_15_out1_ready = branch_15__Buffer_51__ready__0__anchor__in;
	assign branch_15__Buffer_51__ready__0__anchor__out = Buffer_51_in1_ready;
	assign sink_7_in1_data = branch_15__sink_7__data__0__anchor__in;
	assign branch_15__sink_7__data__0__anchor__out = branch_15_out2_data;
	assign sink_7_in1_valid = branch_15__sink_7__valid__0__anchor__in;
	assign branch_15__sink_7__valid__0__anchor__out = branch_15_out2_valid;
	assign branch_15_out2_ready = branch_15__sink_7__ready__0__anchor__in;
	assign branch_15__sink_7__ready__0__anchor__out = sink_7_in1_ready;
	assign branch_16_clk = clk;
	assign branch_16_rst = rst;
	assign Buffer_55_in1_data = branch_16__Buffer_55__data__0__anchor__in;
	assign branch_16__Buffer_55__data__0__anchor__out = branch_16_out1_data;
	assign Buffer_55_in1_valid = branch_16__Buffer_55__valid__0__anchor__in;
	assign branch_16__Buffer_55__valid__0__anchor__out = branch_16_out1_valid;
	assign branch_16_out1_ready = branch_16__Buffer_55__ready__0__anchor__in;
	assign branch_16__Buffer_55__ready__0__anchor__out = Buffer_55_in1_ready;
	assign sink_8_in1_data = branch_16__sink_8__data__0__anchor__in;
	assign branch_16__sink_8__data__0__anchor__out = branch_16_out2_data;
	assign sink_8_in1_valid = branch_16__sink_8__valid__0__anchor__in;
	assign branch_16__sink_8__valid__0__anchor__out = branch_16_out2_valid;
	assign branch_16_out2_ready = branch_16__sink_8__ready__0__anchor__in;
	assign branch_16__sink_8__ready__0__anchor__out = sink_8_in1_ready;
	assign branch_17_clk = clk;
	assign branch_17_rst = rst;
	assign Buffer_54_in1_data = branch_17__Buffer_54__data__0__anchor__in;
	assign branch_17__Buffer_54__data__0__anchor__out = branch_17_out1_data;
	assign Buffer_54_in1_valid = branch_17__Buffer_54__valid__0__anchor__in;
	assign branch_17__Buffer_54__valid__0__anchor__out = branch_17_out1_valid;
	assign branch_17_out1_ready = branch_17__Buffer_54__ready__0__anchor__in;
	assign branch_17__Buffer_54__ready__0__anchor__out = Buffer_54_in1_ready;
	assign sink_9_in1_data = branch_17__sink_9__data__0__anchor__in;
	assign branch_17__sink_9__data__0__anchor__out = branch_17_out2_data;
	assign sink_9_in1_valid = branch_17__sink_9__valid__0__anchor__in;
	assign branch_17__sink_9__valid__0__anchor__out = branch_17_out2_valid;
	assign branch_17_out2_ready = branch_17__sink_9__ready__0__anchor__in;
	assign branch_17__sink_9__ready__0__anchor__out = sink_9_in1_ready;
	assign branch_18_clk = clk;
	assign branch_18_rst = rst;
	assign Buffer_53_in1_data = branch_18__Buffer_53__data__0__anchor__in;
	assign branch_18__Buffer_53__data__0__anchor__out = branch_18_out1_data;
	assign Buffer_53_in1_valid = branch_18__Buffer_53__valid__0__anchor__in;
	assign branch_18__Buffer_53__valid__0__anchor__out = branch_18_out1_valid;
	assign branch_18_out1_ready = branch_18__Buffer_53__ready__0__anchor__in;
	assign branch_18__Buffer_53__ready__0__anchor__out = Buffer_53_in1_ready;
	assign sink_10_in1_data = branch_18__sink_10__data__0__anchor__in;
	assign branch_18__sink_10__data__0__anchor__out = branch_18_out2_data;
	assign sink_10_in1_valid = branch_18__sink_10__valid__0__anchor__in;
	assign branch_18__sink_10__valid__0__anchor__out = branch_18_out2_valid;
	assign branch_18_out2_ready = branch_18__sink_10__ready__0__anchor__in;
	assign branch_18__sink_10__ready__0__anchor__out = sink_10_in1_ready;
	assign fork_18_clk = clk;
	assign fork_18_rst = rst;
	assign branch_18_in2_data = fork_18__branch_18__data__0__anchor__in;
	assign fork_18__branch_18__data__0__anchor__out = fork_18_out1_data;
	assign branch_18_in2_valid = fork_18__branch_18__valid__0__anchor__in;
	assign fork_18__branch_18__valid__0__anchor__out = fork_18_out1_valid;
	assign fork_18_out1_ready = fork_18__branch_18__ready__0__anchor__in;
	assign fork_18__branch_18__ready__0__anchor__out = branch_18_in2_ready;
	assign branch_17_in2_data = fork_18__branch_17__data__0__anchor__in;
	assign fork_18__branch_17__data__0__anchor__out = fork_18_out2_data;
	assign branch_17_in2_valid = fork_18__branch_17__valid__0__anchor__in;
	assign fork_18__branch_17__valid__0__anchor__out = fork_18_out2_valid;
	assign fork_18_out2_ready = fork_18__branch_17__ready__0__anchor__in;
	assign fork_18__branch_17__ready__0__anchor__out = branch_17_in2_ready;
	assign branch_16_in2_data = fork_18__branch_16__data__0__anchor__in;
	assign fork_18__branch_16__data__0__anchor__out = fork_18_out3_data;
	assign branch_16_in2_valid = fork_18__branch_16__valid__0__anchor__in;
	assign fork_18__branch_16__valid__0__anchor__out = fork_18_out3_valid;
	assign fork_18_out3_ready = fork_18__branch_16__ready__0__anchor__in;
	assign fork_18__branch_16__ready__0__anchor__out = branch_16_in2_ready;
	assign branch_15_in2_data = fork_18__branch_15__data__0__anchor__in;
	assign fork_18__branch_15__data__0__anchor__out = fork_18_out4_data;
	assign branch_15_in2_valid = fork_18__branch_15__valid__0__anchor__in;
	assign fork_18__branch_15__valid__0__anchor__out = fork_18_out4_valid;
	assign fork_18_out4_ready = fork_18__branch_15__ready__0__anchor__in;
	assign fork_18__branch_15__ready__0__anchor__out = branch_15_in2_ready;
	assign branchC_26_in2_data = fork_18__branchC_26__data__0__anchor__in;
	assign fork_18__branchC_26__data__0__anchor__out = fork_18_out5_data;
	assign branchC_26_in2_valid = fork_18__branchC_26__valid__0__anchor__in;
	assign fork_18__branchC_26__valid__0__anchor__out = fork_18_out5_valid;
	assign fork_18_out5_ready = fork_18__branchC_26__ready__0__anchor__in;
	assign fork_18__branchC_26__ready__0__anchor__out = branchC_26_in2_ready;
	assign branch_19_clk = clk;
	assign branch_19_rst = rst;
	assign Buffer_52_in1_data = branch_19__Buffer_52__data__0__anchor__in;
	assign branch_19__Buffer_52__data__0__anchor__out = branch_19_out1_data;
	assign Buffer_52_in1_valid = branch_19__Buffer_52__valid__0__anchor__in;
	assign branch_19__Buffer_52__valid__0__anchor__out = branch_19_out1_valid;
	assign branch_19_out1_ready = branch_19__Buffer_52__ready__0__anchor__in;
	assign branch_19__Buffer_52__ready__0__anchor__out = Buffer_52_in1_ready;
	assign sink_11_in1_data = branch_19__sink_11__data__0__anchor__in;
	assign branch_19__sink_11__data__0__anchor__out = branch_19_out2_data;
	assign sink_11_in1_valid = branch_19__sink_11__valid__0__anchor__in;
	assign branch_19__sink_11__valid__0__anchor__out = branch_19_out2_valid;
	assign branch_19_out2_ready = branch_19__sink_11__ready__0__anchor__in;
	assign branch_19__sink_11__ready__0__anchor__out = sink_11_in1_ready;
	assign branch_20_clk = clk;
	assign branch_20_rst = rst;
	assign Buffer_50_in1_data = branch_20__Buffer_50__data__0__anchor__in;
	assign branch_20__Buffer_50__data__0__anchor__out = branch_20_out1_data;
	assign Buffer_50_in1_valid = branch_20__Buffer_50__valid__0__anchor__in;
	assign branch_20__Buffer_50__valid__0__anchor__out = branch_20_out1_valid;
	assign branch_20_out1_ready = branch_20__Buffer_50__ready__0__anchor__in;
	assign branch_20__Buffer_50__ready__0__anchor__out = Buffer_50_in1_ready;
	assign sink_12_in1_data = branch_20__sink_12__data__0__anchor__in;
	assign branch_20__sink_12__data__0__anchor__out = branch_20_out2_data;
	assign sink_12_in1_valid = branch_20__sink_12__valid__0__anchor__in;
	assign branch_20__sink_12__valid__0__anchor__out = branch_20_out2_valid;
	assign branch_20_out2_ready = branch_20__sink_12__ready__0__anchor__in;
	assign branch_20__sink_12__ready__0__anchor__out = sink_12_in1_ready;
	assign fork_19_clk = clk;
	assign fork_19_rst = rst;
	assign branch_20_in2_data = fork_19__branch_20__data__0__anchor__in;
	assign fork_19__branch_20__data__0__anchor__out = fork_19_out1_data;
	assign branch_20_in2_valid = fork_19__branch_20__valid__0__anchor__in;
	assign fork_19__branch_20__valid__0__anchor__out = fork_19_out1_valid;
	assign fork_19_out1_ready = fork_19__branch_20__ready__0__anchor__in;
	assign fork_19__branch_20__ready__0__anchor__out = branch_20_in2_ready;
	assign branch_19_in2_data = fork_19__branch_19__data__0__anchor__in;
	assign fork_19__branch_19__data__0__anchor__out = fork_19_out2_data;
	assign branch_19_in2_valid = fork_19__branch_19__valid__0__anchor__in;
	assign fork_19__branch_19__valid__0__anchor__out = fork_19_out2_valid;
	assign fork_19_out2_ready = fork_19__branch_19__ready__0__anchor__in;
	assign fork_19__branch_19__ready__0__anchor__out = branch_19_in2_ready;
	assign branchC_27_in2_data = fork_19__branchC_27__data__0__anchor__in;
	assign fork_19__branchC_27__data__0__anchor__out = fork_19_out3_data;
	assign branchC_27_in2_valid = fork_19__branchC_27__valid__0__anchor__in;
	assign fork_19__branchC_27__valid__0__anchor__out = fork_19_out3_valid;
	assign fork_19_out3_ready = fork_19__branchC_27__ready__0__anchor__in;
	assign fork_19__branchC_27__ready__0__anchor__out = branchC_27_in2_ready;
	assign MC_A_clk = clk;
	assign MC_A_rst = rst;
	assign A_ce0 = A_we0;
	assign load_6_in1_data = MC_A__load_6__data__0__anchor__in;
	assign MC_A__load_6__data__0__anchor__out = MC_A_out1_data;
	assign load_6_in1_valid = MC_A__load_6__valid__0__anchor__in;
	assign MC_A__load_6__valid__0__anchor__out = MC_A_out1_valid;
	assign MC_A_out1_ready = MC_A__load_6__ready__0__anchor__in;
	assign MC_A__load_6__ready__0__anchor__out = load_6_in1_ready;
	assign load_14_in1_data = MC_A__load_14__data__0__anchor__in;
	assign MC_A__load_14__data__0__anchor__out = MC_A_out2_data;
	assign load_14_in1_valid = MC_A__load_14__valid__0__anchor__in;
	assign MC_A__load_14__valid__0__anchor__out = MC_A_out2_valid;
	assign MC_A_out2_ready = MC_A__load_14__ready__0__anchor__in;
	assign MC_A__load_14__ready__0__anchor__out = load_14_in1_ready;
	assign load_20_in1_data = MC_A__load_20__data__0__anchor__in;
	assign MC_A__load_20__data__0__anchor__out = MC_A_out3_data;
	assign load_20_in1_valid = MC_A__load_20__valid__0__anchor__in;
	assign MC_A__load_20__valid__0__anchor__out = MC_A_out3_valid;
	assign MC_A_out3_ready = MC_A__load_20__ready__0__anchor__in;
	assign MC_A__load_20__ready__0__anchor__out = load_20_in1_ready;
	assign end_0_in1_data = MC_A__end_0__data__0__anchor__in;
	assign MC_A__end_0__data__0__anchor__out = MC_A_out4_data;
	assign end_0_in1_valid = MC_A__end_0__valid__0__anchor__in;
	assign MC_A__end_0__valid__0__anchor__out = MC_A_out4_valid;
	assign MC_A_out4_ready = MC_A__end_0__ready__0__anchor__in;
	assign MC_A__end_0__ready__0__anchor__out = end_0_in1_ready;
	assign cst_7_clk = clk;
	assign cst_7_rst = rst;
	assign MC_A_in1_data = cst_7__MC_A__data__0__anchor__in;
	assign cst_7__MC_A__data__0__anchor__out = cst_7_out1_data;
	assign MC_A_in1_valid = cst_7__MC_A__valid__0__anchor__in;
	assign cst_7__MC_A__valid__0__anchor__out = cst_7_out1_valid;
	assign cst_7_out1_ready = cst_7__MC_A__ready__0__anchor__in;
	assign cst_7__MC_A__ready__0__anchor__out = MC_A_in1_ready;
	assign cst_8_clk = clk;
	assign cst_8_rst = rst;
	assign MC_A_in2_data = cst_8__MC_A__data__0__anchor__in;
	assign cst_8__MC_A__data__0__anchor__out = cst_8_out1_data;
	assign MC_A_in2_valid = cst_8__MC_A__valid__0__anchor__in;
	assign cst_8__MC_A__valid__0__anchor__out = cst_8_out1_valid;
	assign cst_8_out1_ready = cst_8__MC_A__ready__0__anchor__in;
	assign cst_8__MC_A__ready__0__anchor__out = MC_A_in2_ready;
	assign end_0_clk = clk;
	assign end_0_rst = rst;
	assign end_out = end_0_out1_data;
	assign end_0_out1_ready = end_ready;
	assign end_valid = end_0_out1_valid;
	assign start_0_clk = clk;
	assign start_0_rst = rst;
	assign start_0_in1_data = start_in;
	assign start_0_in1_valid = start_valid;
	assign start_ready = start_0_in1_ready;
	assign branchC_21_in1_data = start_0__branchC_21__data__0__anchor__in;
	assign start_0__branchC_21__data__0__anchor__out = start_0_out1_data;
	assign branchC_21_in1_valid = start_0__branchC_21__valid__0__anchor__in;
	assign start_0__branchC_21__valid__0__anchor__out = start_0_out1_valid;
	assign start_0_out1_ready = start_0__branchC_21__ready__0__anchor__in;
	assign start_0__branchC_21__ready__0__anchor__out = branchC_21_in1_ready;
	assign branchC_21_clk = clk;
	assign branchC_21_rst = rst;
	assign phiC_23_in1_data = branchC_21__phiC_23__data__0__anchor__in;
	assign branchC_21__phiC_23__data__0__anchor__out = branchC_21_out1_data;
	assign phiC_23_in1_valid = branchC_21__phiC_23__valid__0__anchor__in;
	assign branchC_21__phiC_23__valid__0__anchor__out = branchC_21_out1_valid;
	assign branchC_21_out1_ready = branchC_21__phiC_23__ready__0__anchor__in;
	assign branchC_21__phiC_23__ready__0__anchor__out = phiC_23_in1_ready;
	assign phiC_17_in1_data = branchC_21__phiC_17__data__0__anchor__in;
	assign branchC_21__phiC_17__data__0__anchor__out = branchC_21_out2_data;
	assign phiC_17_in1_valid = branchC_21__phiC_17__valid__0__anchor__in;
	assign branchC_21__phiC_17__valid__0__anchor__out = branchC_21_out2_valid;
	assign branchC_21_out2_ready = branchC_21__phiC_17__ready__0__anchor__in;
	assign branchC_21__phiC_17__ready__0__anchor__out = phiC_17_in1_ready;
	assign fork_22_clk = clk;
	assign fork_22_rst = rst;
	assign branch_0_in2_data = fork_22__branch_0__data__0__anchor__in;
	assign fork_22__branch_0__data__0__anchor__out = fork_22_out1_data;
	assign branch_0_in2_valid = fork_22__branch_0__valid__0__anchor__in;
	assign fork_22__branch_0__valid__0__anchor__out = fork_22_out1_valid;
	assign fork_22_out1_ready = fork_22__branch_0__ready__0__anchor__in;
	assign fork_22__branch_0__ready__0__anchor__out = branch_0_in2_ready;
	assign branchC_21_in2_data = fork_22__branchC_21__data__0__anchor__in;
	assign fork_22__branchC_21__data__0__anchor__out = fork_22_out2_data;
	assign branchC_21_in2_valid = fork_22__branchC_21__valid__0__anchor__in;
	assign fork_22__branchC_21__valid__0__anchor__out = fork_22_out2_valid;
	assign fork_22_out2_ready = fork_22__branchC_21__ready__0__anchor__in;
	assign fork_22__branchC_21__ready__0__anchor__out = branchC_21_in2_ready;
	assign phiC_17_clk = clk;
	assign phiC_17_rst = rst;
	assign forkC_23_in1_data = phiC_17__forkC_23__data__0__anchor__in;
	assign phiC_17__forkC_23__data__0__anchor__out = phiC_17_out1_data;
	assign forkC_23_in1_valid = phiC_17__forkC_23__valid__0__anchor__in;
	assign phiC_17__forkC_23__valid__0__anchor__out = phiC_17_out1_valid;
	assign phiC_17_out1_ready = phiC_17__forkC_23__ready__0__anchor__in;
	assign phiC_17__forkC_23__ready__0__anchor__out = forkC_23_in1_ready;
	assign forkC_23_clk = clk;
	assign forkC_23_rst = rst;
	assign cst_1_in1_data = forkC_23__cst_1__data__0__anchor__in;
	assign forkC_23__cst_1__data__0__anchor__out = forkC_23_out1_data;
	assign cst_1_in1_valid = forkC_23__cst_1__valid__0__anchor__in;
	assign forkC_23__cst_1__valid__0__anchor__out = forkC_23_out1_valid;
	assign forkC_23_out1_ready = forkC_23__cst_1__ready__0__anchor__in;
	assign forkC_23__cst_1__ready__0__anchor__out = cst_1_in1_ready;
	assign branchC_22_in1_data = forkC_23__branchC_22__data__0__anchor__in;
	assign forkC_23__branchC_22__data__0__anchor__out = forkC_23_out2_data;
	assign branchC_22_in1_valid = forkC_23__branchC_22__valid__0__anchor__in;
	assign forkC_23__branchC_22__valid__0__anchor__out = forkC_23_out2_valid;
	assign forkC_23_out2_ready = forkC_23__branchC_22__ready__0__anchor__in;
	assign forkC_23__branchC_22__ready__0__anchor__out = branchC_22_in1_ready;
	assign brCst_block2_in1_data = forkC_23__brCst_block2__data__0__anchor__in;
	assign forkC_23__brCst_block2__data__0__anchor__out = forkC_23_out3_data;
	assign brCst_block2_in1_valid = forkC_23__brCst_block2__valid__0__anchor__in;
	assign forkC_23__brCst_block2__valid__0__anchor__out = forkC_23_out3_valid;
	assign forkC_23_out3_ready = forkC_23__brCst_block2__ready__0__anchor__in;
	assign forkC_23__brCst_block2__ready__0__anchor__out = brCst_block2_in1_ready;
	assign branchC_22_clk = clk;
	assign branchC_22_rst = rst;
	assign phiC_18_in1_data = branchC_22__phiC_18__data__0__anchor__in;
	assign branchC_22__phiC_18__data__0__anchor__out = branchC_22_out1_data;
	assign phiC_18_in1_valid = branchC_22__phiC_18__valid__0__anchor__in;
	assign branchC_22__phiC_18__valid__0__anchor__out = branchC_22_out1_valid;
	assign branchC_22_out1_ready = branchC_22__phiC_18__ready__0__anchor__in;
	assign branchC_22__phiC_18__ready__0__anchor__out = phiC_18_in1_ready;
	assign sink_13_in1_data = branchC_22__sink_13__data__0__anchor__in;
	assign branchC_22__sink_13__data__0__anchor__out = branchC_22_out2_data;
	assign sink_13_in1_valid = branchC_22__sink_13__valid__0__anchor__in;
	assign branchC_22__sink_13__valid__0__anchor__out = branchC_22_out2_valid;
	assign branchC_22_out2_ready = branchC_22__sink_13__ready__0__anchor__in;
	assign branchC_22__sink_13__ready__0__anchor__out = sink_13_in1_ready;
	assign phiC_18_clk = clk;
	assign phiC_18_rst = rst;
	assign forkC_24_in1_data = phiC_18__forkC_24__data__0__anchor__in;
	assign phiC_18__forkC_24__data__0__anchor__out = phiC_18_out1_data;
	assign forkC_24_in1_valid = phiC_18__forkC_24__valid__0__anchor__in;
	assign phiC_18__forkC_24__valid__0__anchor__out = phiC_18_out1_valid;
	assign phiC_18_out1_ready = phiC_18__forkC_24__ready__0__anchor__in;
	assign phiC_18__forkC_24__ready__0__anchor__out = forkC_24_in1_ready;
	assign phi_3_in1_data = phiC_18__phi_3__data__0__anchor__in;
	assign phiC_18__phi_3__data__0__anchor__out = phiC_18_out2_data;
	assign phi_3_in1_valid = phiC_18__phi_3__valid__0__anchor__in;
	assign phiC_18__phi_3__valid__0__anchor__out = phiC_18_out2_valid;
	assign phiC_18_out2_ready = phiC_18__phi_3__ready__0__anchor__in;
	assign phiC_18__phi_3__ready__0__anchor__out = phi_3_in1_ready;
	assign forkC_24_clk = clk;
	assign forkC_24_rst = rst;
	assign branchC_23_in1_data = forkC_24__branchC_23__data__0__anchor__in;
	assign forkC_24__branchC_23__data__0__anchor__out = forkC_24_out1_data;
	assign branchC_23_in1_valid = forkC_24__branchC_23__valid__0__anchor__in;
	assign forkC_24__branchC_23__valid__0__anchor__out = forkC_24_out1_valid;
	assign forkC_24_out1_ready = forkC_24__branchC_23__ready__0__anchor__in;
	assign forkC_24__branchC_23__ready__0__anchor__out = branchC_23_in1_ready;
	assign brCst_block3_in1_data = forkC_24__brCst_block3__data__0__anchor__in;
	assign forkC_24__brCst_block3__data__0__anchor__out = forkC_24_out2_data;
	assign brCst_block3_in1_valid = forkC_24__brCst_block3__valid__0__anchor__in;
	assign forkC_24__brCst_block3__valid__0__anchor__out = forkC_24_out2_valid;
	assign forkC_24_out2_ready = forkC_24__brCst_block3__ready__0__anchor__in;
	assign forkC_24__brCst_block3__ready__0__anchor__out = brCst_block3_in1_ready;
	assign branchC_23_clk = clk;
	assign branchC_23_rst = rst;
	assign phiC_19_in1_data = branchC_23__phiC_19__data__0__anchor__in;
	assign branchC_23__phiC_19__data__0__anchor__out = branchC_23_out1_data;
	assign phiC_19_in1_valid = branchC_23__phiC_19__valid__0__anchor__in;
	assign branchC_23__phiC_19__valid__0__anchor__out = branchC_23_out1_valid;
	assign branchC_23_out1_ready = branchC_23__phiC_19__ready__0__anchor__in;
	assign branchC_23__phiC_19__ready__0__anchor__out = phiC_19_in1_ready;
	assign sink_14_in1_data = branchC_23__sink_14__data__0__anchor__in;
	assign branchC_23__sink_14__data__0__anchor__out = branchC_23_out2_data;
	assign sink_14_in1_valid = branchC_23__sink_14__valid__0__anchor__in;
	assign branchC_23__sink_14__valid__0__anchor__out = branchC_23_out2_valid;
	assign branchC_23_out2_ready = branchC_23__sink_14__ready__0__anchor__in;
	assign branchC_23__sink_14__ready__0__anchor__out = sink_14_in1_ready;
	assign phiC_19_clk = clk;
	assign phiC_19_rst = rst;
	assign branchC_24_in1_data = phiC_19__branchC_24__data__0__anchor__in;
	assign phiC_19__branchC_24__data__0__anchor__out = phiC_19_out1_data;
	assign branchC_24_in1_valid = phiC_19__branchC_24__valid__0__anchor__in;
	assign phiC_19__branchC_24__valid__0__anchor__out = phiC_19_out1_valid;
	assign phiC_19_out1_ready = phiC_19__branchC_24__ready__0__anchor__in;
	assign phiC_19__branchC_24__ready__0__anchor__out = branchC_24_in1_ready;
	assign phi_8_in1_data = phiC_19__phi_8__data__0__anchor__in;
	assign phiC_19__phi_8__data__0__anchor__out = phiC_19_out2_data;
	assign phi_8_in1_valid = phiC_19__phi_8__valid__0__anchor__in;
	assign phiC_19__phi_8__valid__0__anchor__out = phiC_19_out2_valid;
	assign phiC_19_out2_ready = phiC_19__phi_8__ready__0__anchor__in;
	assign phiC_19__phi_8__ready__0__anchor__out = phi_8_in1_ready;
	assign branchC_24_clk = clk;
	assign branchC_24_rst = rst;
	assign phiC_20_in1_data = branchC_24__phiC_20__data__0__anchor__in;
	assign branchC_24__phiC_20__data__0__anchor__out = branchC_24_out1_data;
	assign phiC_20_in1_valid = branchC_24__phiC_20__valid__0__anchor__in;
	assign branchC_24__phiC_20__valid__0__anchor__out = branchC_24_out1_valid;
	assign branchC_24_out1_ready = branchC_24__phiC_20__ready__0__anchor__in;
	assign branchC_24__phiC_20__ready__0__anchor__out = phiC_20_in1_ready;
	assign phiC_22_in1_data = branchC_24__phiC_22__data__0__anchor__in;
	assign branchC_24__phiC_22__data__0__anchor__out = branchC_24_out2_data;
	assign phiC_22_in1_valid = branchC_24__phiC_22__valid__0__anchor__in;
	assign branchC_24__phiC_22__valid__0__anchor__out = branchC_24_out2_valid;
	assign branchC_24_out2_ready = branchC_24__phiC_22__ready__0__anchor__in;
	assign branchC_24__phiC_22__ready__0__anchor__out = phiC_22_in1_ready;
	assign phiC_20_clk = clk;
	assign phiC_20_rst = rst;
	assign branchC_25_in1_data = phiC_20__branchC_25__data__0__anchor__in;
	assign phiC_20__branchC_25__data__0__anchor__out = phiC_20_out1_data;
	assign branchC_25_in1_valid = phiC_20__branchC_25__valid__0__anchor__in;
	assign phiC_20__branchC_25__valid__0__anchor__out = phiC_20_out1_valid;
	assign phiC_20_out1_ready = phiC_20__branchC_25__ready__0__anchor__in;
	assign phiC_20__branchC_25__ready__0__anchor__out = branchC_25_in1_ready;
	assign branchC_25_clk = clk;
	assign branchC_25_rst = rst;
	assign phiC_21_in1_data = branchC_25__phiC_21__data__0__anchor__in;
	assign branchC_25__phiC_21__data__0__anchor__out = branchC_25_out1_data;
	assign phiC_21_in1_valid = branchC_25__phiC_21__valid__0__anchor__in;
	assign branchC_25__phiC_21__valid__0__anchor__out = branchC_25_out1_valid;
	assign branchC_25_out1_ready = branchC_25__phiC_21__ready__0__anchor__in;
	assign branchC_25__phiC_21__ready__0__anchor__out = phiC_21_in1_ready;
	assign phiC_22_in2_data = branchC_25__phiC_22__data__0__anchor__in;
	assign branchC_25__phiC_22__data__0__anchor__out = branchC_25_out2_data;
	assign phiC_22_in2_valid = branchC_25__phiC_22__valid__0__anchor__in;
	assign branchC_25__phiC_22__valid__0__anchor__out = branchC_25_out2_valid;
	assign branchC_25_out2_ready = branchC_25__phiC_22__ready__0__anchor__in;
	assign branchC_25__phiC_22__ready__0__anchor__out = phiC_22_in2_ready;
	assign phiC_21_clk = clk;
	assign phiC_21_rst = rst;
	assign forkC_27_in1_data = phiC_21__forkC_27__data__0__anchor__in;
	assign phiC_21__forkC_27__data__0__anchor__out = phiC_21_out1_data;
	assign forkC_27_in1_valid = phiC_21__forkC_27__valid__0__anchor__in;
	assign phiC_21__forkC_27__valid__0__anchor__out = phiC_21_out1_valid;
	assign phiC_21_out1_ready = phiC_21__forkC_27__ready__0__anchor__in;
	assign phiC_21__forkC_27__ready__0__anchor__out = forkC_27_in1_ready;
	assign forkC_27_clk = clk;
	assign forkC_27_rst = rst;
	assign cst_7_in1_data = forkC_27__cst_7__data__0__anchor__in;
	assign forkC_27__cst_7__data__0__anchor__out = forkC_27_out1_data;
	assign cst_7_in1_valid = forkC_27__cst_7__valid__0__anchor__in;
	assign forkC_27__cst_7__valid__0__anchor__out = forkC_27_out1_valid;
	assign forkC_27_out1_ready = forkC_27__cst_7__ready__0__anchor__in;
	assign forkC_27__cst_7__ready__0__anchor__out = cst_7_in1_ready;
	assign branchC_26_in1_data = forkC_27__branchC_26__data__0__anchor__in;
	assign forkC_27__branchC_26__data__0__anchor__out = forkC_27_out2_data;
	assign branchC_26_in1_valid = forkC_27__branchC_26__valid__0__anchor__in;
	assign forkC_27__branchC_26__valid__0__anchor__out = forkC_27_out2_valid;
	assign forkC_27_out2_ready = forkC_27__branchC_26__ready__0__anchor__in;
	assign forkC_27__branchC_26__ready__0__anchor__out = branchC_26_in1_ready;
	assign brCst_block6_in1_data = forkC_27__brCst_block6__data__0__anchor__in;
	assign forkC_27__brCst_block6__data__0__anchor__out = forkC_27_out3_data;
	assign brCst_block6_in1_valid = forkC_27__brCst_block6__valid__0__anchor__in;
	assign forkC_27__brCst_block6__valid__0__anchor__out = forkC_27_out3_valid;
	assign forkC_27_out3_ready = forkC_27__brCst_block6__ready__0__anchor__in;
	assign forkC_27__brCst_block6__ready__0__anchor__out = brCst_block6_in1_ready;
	assign branchC_26_clk = clk;
	assign branchC_26_rst = rst;
	assign Buffer_57_in1_data = branchC_26__Buffer_57__data__0__anchor__in;
	assign branchC_26__Buffer_57__data__0__anchor__out = branchC_26_out1_data;
	assign Buffer_57_in1_valid = branchC_26__Buffer_57__valid__0__anchor__in;
	assign branchC_26__Buffer_57__valid__0__anchor__out = branchC_26_out1_valid;
	assign branchC_26_out1_ready = branchC_26__Buffer_57__ready__0__anchor__in;
	assign branchC_26__Buffer_57__ready__0__anchor__out = Buffer_57_in1_ready;
	assign sink_15_in1_data = branchC_26__sink_15__data__0__anchor__in;
	assign branchC_26__sink_15__data__0__anchor__out = branchC_26_out2_data;
	assign sink_15_in1_valid = branchC_26__sink_15__valid__0__anchor__in;
	assign branchC_26__sink_15__valid__0__anchor__out = branchC_26_out2_valid;
	assign branchC_26_out2_ready = branchC_26__sink_15__ready__0__anchor__in;
	assign branchC_26__sink_15__ready__0__anchor__out = sink_15_in1_ready;
	assign phiC_22_clk = clk;
	assign phiC_22_rst = rst;
	assign forkC_28_in1_data = phiC_22__forkC_28__data__0__anchor__in;
	assign phiC_22__forkC_28__data__0__anchor__out = phiC_22_out1_data;
	assign forkC_28_in1_valid = phiC_22__forkC_28__valid__0__anchor__in;
	assign phiC_22__forkC_28__valid__0__anchor__out = phiC_22_out1_valid;
	assign phiC_22_out1_ready = phiC_22__forkC_28__ready__0__anchor__in;
	assign phiC_22__forkC_28__ready__0__anchor__out = forkC_28_in1_ready;
	assign forkC_28_clk = clk;
	assign forkC_28_rst = rst;
	assign cst_8_in1_data = forkC_28__cst_8__data__0__anchor__in;
	assign forkC_28__cst_8__data__0__anchor__out = forkC_28_out1_data;
	assign cst_8_in1_valid = forkC_28__cst_8__valid__0__anchor__in;
	assign forkC_28__cst_8__valid__0__anchor__out = forkC_28_out1_valid;
	assign forkC_28_out1_ready = forkC_28__cst_8__ready__0__anchor__in;
	assign forkC_28__cst_8__ready__0__anchor__out = cst_8_in1_ready;
	assign branchC_27_in1_data = forkC_28__branchC_27__data__0__anchor__in;
	assign forkC_28__branchC_27__data__0__anchor__out = forkC_28_out2_data;
	assign branchC_27_in1_valid = forkC_28__branchC_27__valid__0__anchor__in;
	assign forkC_28__branchC_27__valid__0__anchor__out = forkC_28_out2_valid;
	assign forkC_28_out2_ready = forkC_28__branchC_27__ready__0__anchor__in;
	assign forkC_28__branchC_27__ready__0__anchor__out = branchC_27_in1_ready;
	assign branchC_27_clk = clk;
	assign branchC_27_rst = rst;
	assign Buffer_56_in1_data = branchC_27__Buffer_56__data__0__anchor__in;
	assign branchC_27__Buffer_56__data__0__anchor__out = branchC_27_out1_data;
	assign Buffer_56_in1_valid = branchC_27__Buffer_56__valid__0__anchor__in;
	assign branchC_27__Buffer_56__valid__0__anchor__out = branchC_27_out1_valid;
	assign branchC_27_out1_ready = branchC_27__Buffer_56__ready__0__anchor__in;
	assign branchC_27__Buffer_56__ready__0__anchor__out = Buffer_56_in1_ready;
	assign phiC_23_in2_data = branchC_27__phiC_23__data__0__anchor__in;
	assign branchC_27__phiC_23__data__0__anchor__out = branchC_27_out2_data;
	assign phiC_23_in2_valid = branchC_27__phiC_23__valid__0__anchor__in;
	assign branchC_27__phiC_23__valid__0__anchor__out = branchC_27_out2_valid;
	assign branchC_27_out2_ready = branchC_27__phiC_23__ready__0__anchor__in;
	assign branchC_27__phiC_23__ready__0__anchor__out = phiC_23_in2_ready;
	assign phiC_23_clk = clk;
	assign phiC_23_rst = rst;
	assign ret_0_in1_data = phiC_23__ret_0__data__0__anchor__in;
	assign phiC_23__ret_0__data__0__anchor__out = phiC_23_out1_data;
	assign ret_0_in1_valid = phiC_23__ret_0__valid__0__anchor__in;
	assign phiC_23__ret_0__valid__0__anchor__out = phiC_23_out1_valid;
	assign phiC_23_out1_ready = phiC_23__ret_0__ready__0__anchor__in;
	assign phiC_23__ret_0__ready__0__anchor__out = ret_0_in1_ready;
	assign sink_0_clk = clk;
	assign sink_0_rst = rst;
	assign sink_1_clk = clk;
	assign sink_1_rst = rst;
	assign sink_2_clk = clk;
	assign sink_2_rst = rst;
	assign sink_3_clk = clk;
	assign sink_3_rst = rst;
	assign sink_4_clk = clk;
	assign sink_4_rst = rst;
	assign sink_5_clk = clk;
	assign sink_5_rst = rst;
	assign sink_6_clk = clk;
	assign sink_6_rst = rst;
	assign sink_7_clk = clk;
	assign sink_7_rst = rst;
	assign sink_8_clk = clk;
	assign sink_8_rst = rst;
	assign sink_9_clk = clk;
	assign sink_9_rst = rst;
	assign sink_10_clk = clk;
	assign sink_10_rst = rst;
	assign sink_11_clk = clk;
	assign sink_11_rst = rst;
	assign sink_12_clk = clk;
	assign sink_12_rst = rst;
	assign sink_13_clk = clk;
	assign sink_13_rst = rst;
	assign sink_14_clk = clk;
	assign sink_14_rst = rst;
	assign sink_15_clk = clk;
	assign sink_15_rst = rst;
	assign source_0_clk = clk;
	assign source_0_rst = rst;
	assign cst_0_in1_data = source_0__cst_0__data__0__anchor__in;
	assign source_0__cst_0__data__0__anchor__out = source_0_out1_data;
	assign cst_0_in1_valid = source_0__cst_0__valid__0__anchor__in;
	assign source_0__cst_0__valid__0__anchor__out = source_0_out1_valid;
	assign source_0_out1_ready = source_0__cst_0__ready__0__anchor__in;
	assign source_0__cst_0__ready__0__anchor__out = cst_0_in1_ready;
	assign source_1_clk = clk;
	assign source_1_rst = rst;
	assign cst_2_in1_data = source_1__cst_2__data__0__anchor__in;
	assign source_1__cst_2__data__0__anchor__out = source_1_out1_data;
	assign cst_2_in1_valid = source_1__cst_2__valid__0__anchor__in;
	assign source_1__cst_2__valid__0__anchor__out = source_1_out1_valid;
	assign source_1_out1_ready = source_1__cst_2__ready__0__anchor__in;
	assign source_1__cst_2__ready__0__anchor__out = cst_2_in1_ready;
	assign source_2_clk = clk;
	assign source_2_rst = rst;
	assign cst_3_in1_data = source_2__cst_3__data__0__anchor__in;
	assign source_2__cst_3__data__0__anchor__out = source_2_out1_data;
	assign cst_3_in1_valid = source_2__cst_3__valid__0__anchor__in;
	assign source_2__cst_3__valid__0__anchor__out = source_2_out1_valid;
	assign source_2_out1_ready = source_2__cst_3__ready__0__anchor__in;
	assign source_2__cst_3__ready__0__anchor__out = cst_3_in1_ready;
	assign source_3_clk = clk;
	assign source_3_rst = rst;
	assign cst_4_in1_data = source_3__cst_4__data__0__anchor__in;
	assign source_3__cst_4__data__0__anchor__out = source_3_out1_data;
	assign cst_4_in1_valid = source_3__cst_4__valid__0__anchor__in;
	assign source_3__cst_4__valid__0__anchor__out = source_3_out1_valid;
	assign source_3_out1_ready = source_3__cst_4__ready__0__anchor__in;
	assign source_3__cst_4__ready__0__anchor__out = cst_4_in1_ready;
	assign source_4_clk = clk;
	assign source_4_rst = rst;
	assign cst_5_in1_data = source_4__cst_5__data__0__anchor__in;
	assign source_4__cst_5__data__0__anchor__out = source_4_out1_data;
	assign cst_5_in1_valid = source_4__cst_5__valid__0__anchor__in;
	assign source_4__cst_5__valid__0__anchor__out = source_4_out1_valid;
	assign source_4_out1_ready = source_4__cst_5__ready__0__anchor__in;
	assign source_4__cst_5__ready__0__anchor__out = cst_5_in1_ready;
	assign source_5_clk = clk;
	assign source_5_rst = rst;
	assign cst_6_in1_data = source_5__cst_6__data__0__anchor__in;
	assign source_5__cst_6__data__0__anchor__out = source_5_out1_data;
	assign cst_6_in1_valid = source_5__cst_6__valid__0__anchor__in;
	assign source_5__cst_6__valid__0__anchor__out = source_5_out1_valid;
	assign source_5_out1_ready = source_5__cst_6__ready__0__anchor__in;
	assign source_5__cst_6__ready__0__anchor__out = cst_6_in1_ready;
	assign Buffer_50_clk = clk;
	assign Buffer_50_rst = rst;
	assign phi_n1_in2_data = Buffer_50__phi_n1__data__0__anchor__in;
	assign Buffer_50__phi_n1__data__0__anchor__out = Buffer_50_out1_data;
	assign phi_n1_in2_valid = Buffer_50__phi_n1__valid__0__anchor__in;
	assign Buffer_50__phi_n1__valid__0__anchor__out = Buffer_50_out1_valid;
	assign Buffer_50_out1_ready = Buffer_50__phi_n1__ready__0__anchor__in;
	assign Buffer_50__phi_n1__ready__0__anchor__out = phi_n1_in2_ready;
	assign Buffer_51_clk = clk;
	assign Buffer_51_rst = rst;
	assign phi_8_in3_data = Buffer_51__phi_8__data__0__anchor__in;
	assign Buffer_51__phi_8__data__0__anchor__out = Buffer_51_out1_data;
	assign phi_8_in3_valid = Buffer_51__phi_8__valid__0__anchor__in;
	assign Buffer_51__phi_8__valid__0__anchor__out = Buffer_51_out1_valid;
	assign Buffer_51_out1_ready = Buffer_51__phi_8__ready__0__anchor__in;
	assign Buffer_51__phi_8__ready__0__anchor__out = phi_8_in3_ready;
	assign Buffer_52_clk = clk;
	assign Buffer_52_rst = rst;
	assign phi_3_in3_data = Buffer_52__phi_3__data__0__anchor__in;
	assign Buffer_52__phi_3__data__0__anchor__out = Buffer_52_out1_data;
	assign phi_3_in3_valid = Buffer_52__phi_3__valid__0__anchor__in;
	assign Buffer_52__phi_3__valid__0__anchor__out = Buffer_52_out1_valid;
	assign Buffer_52_out1_ready = Buffer_52__phi_3__ready__0__anchor__in;
	assign Buffer_52__phi_3__ready__0__anchor__out = phi_3_in3_ready;
	assign Buffer_53_clk = clk;
	assign Buffer_53_rst = rst;
	assign phi_n8_in2_data = Buffer_53__phi_n8__data__0__anchor__in;
	assign Buffer_53__phi_n8__data__0__anchor__out = Buffer_53_out1_data;
	assign phi_n8_in2_valid = Buffer_53__phi_n8__valid__0__anchor__in;
	assign Buffer_53__phi_n8__valid__0__anchor__out = Buffer_53_out1_valid;
	assign Buffer_53_out1_ready = Buffer_53__phi_n8__ready__0__anchor__in;
	assign Buffer_53__phi_n8__ready__0__anchor__out = phi_n8_in2_ready;
	assign Buffer_54_clk = clk;
	assign Buffer_54_rst = rst;
	assign phi_n7_in2_data = Buffer_54__phi_n7__data__0__anchor__in;
	assign Buffer_54__phi_n7__data__0__anchor__out = Buffer_54_out1_data;
	assign phi_n7_in2_valid = Buffer_54__phi_n7__valid__0__anchor__in;
	assign Buffer_54__phi_n7__valid__0__anchor__out = Buffer_54_out1_valid;
	assign Buffer_54_out1_ready = Buffer_54__phi_n7__ready__0__anchor__in;
	assign Buffer_54__phi_n7__ready__0__anchor__out = phi_n7_in2_ready;
	assign Buffer_55_clk = clk;
	assign Buffer_55_rst = rst;
	assign phi_n6_in2_data = Buffer_55__phi_n6__data__0__anchor__in;
	assign Buffer_55__phi_n6__data__0__anchor__out = Buffer_55_out1_data;
	assign phi_n6_in2_valid = Buffer_55__phi_n6__valid__0__anchor__in;
	assign Buffer_55__phi_n6__valid__0__anchor__out = Buffer_55_out1_valid;
	assign Buffer_55_out1_ready = Buffer_55__phi_n6__ready__0__anchor__in;
	assign Buffer_55__phi_n6__ready__0__anchor__out = phi_n6_in2_ready;
	assign Buffer_56_clk = clk;
	assign Buffer_56_rst = rst;
	assign phiC_18_in2_data = Buffer_56__phiC_18__data__0__anchor__in;
	assign Buffer_56__phiC_18__data__0__anchor__out = Buffer_56_out1_data;
	assign phiC_18_in2_valid = Buffer_56__phiC_18__valid__0__anchor__in;
	assign Buffer_56__phiC_18__valid__0__anchor__out = Buffer_56_out1_valid;
	assign Buffer_56_out1_ready = Buffer_56__phiC_18__ready__0__anchor__in;
	assign Buffer_56__phiC_18__ready__0__anchor__out = phiC_18_in2_ready;
	assign Buffer_57_clk = clk;
	assign Buffer_57_rst = rst;
	assign phiC_19_in2_data = Buffer_57__phiC_19__data__0__anchor__in;
	assign Buffer_57__phiC_19__data__0__anchor__out = Buffer_57_out1_data;
	assign phiC_19_in2_valid = Buffer_57__phiC_19__valid__0__anchor__in;
	assign Buffer_57__phiC_19__valid__0__anchor__out = Buffer_57_out1_valid;
	assign Buffer_57_out1_ready = Buffer_57__phiC_19__ready__0__anchor__in;
	assign Buffer_57__phiC_19__ready__0__anchor__out = phiC_19_in2_ready;
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_17 (.clk(phiC_17_clk), .rst(phiC_17_rst), .data_in_bus({phiC_17_in1_data}), .valid_in_bus({phiC_17_in1_valid}), .ready_in_bus({phiC_17_in1_ready}), .data_out_bus({phiC_17_out1_data}), .valid_out_bus({phiC_17_out1_valid}), .ready_out_bus({phiC_17_out1_ready}));
MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(32), .BB_COUNT(2), .LOAD_COUNT(3), .STORE_COUNT(2))MemCont_MC_A (.clk(MC_A_clk), .rst(MC_A_rst), .io_storeDataOut(A_dout0), .io_storeAddrOut(A_address0), .io_storeEnable(A_we0), .io_loadDataIn(A_din1), .io_loadAddrOut(A_address1), .io_loadEnable(A_ce1), .io_bbpValids({MC_A_in2_valid, MC_A_in1_valid}), .io_bb_stCountArray({MC_A_in2_data, MC_A_in1_data}), .io_bbReadyToPrevs({MC_A_in2_ready, MC_A_in1_ready}), .io_rdPortsPrev_ready({MC_A_in5_ready, MC_A_in4_ready, MC_A_in3_ready}), .io_rdPortsPrev_valid({MC_A_in5_valid, MC_A_in4_valid, MC_A_in3_valid}), .io_rdPortsPrev_bits({MC_A_in5_data, MC_A_in4_data, MC_A_in3_data}), .io_wrAddrPorts_ready({MC_A_in8_ready, MC_A_in6_ready}), .io_wrAddrPorts_valid({MC_A_in8_valid, MC_A_in6_valid}), .io_wrAddrPorts_bits({MC_A_in8_data, MC_A_in6_data}), .io_wrDataPorts_ready({MC_A_in9_ready, MC_A_in7_ready}), .io_wrDataPorts_valid({MC_A_in9_valid, MC_A_in7_valid}), .io_wrDataPorts_bits({MC_A_in9_data, MC_A_in7_data}), .io_rdPortsNext_ready({MC_A_out3_ready, MC_A_out2_ready, MC_A_out1_ready}), .io_rdPortsNext_valid({MC_A_out3_valid, MC_A_out2_valid, MC_A_out1_valid}), .io_rdPortsNext_bits({MC_A_out3_data, MC_A_out2_data, MC_A_out1_data}), .io_Empty_Valid({MC_A_out4_valid}), .io_Empty_Ready({MC_A_out4_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_18 (.clk(branch_18_clk), .rst(branch_18_rst), .data_in_bus({{31'b0, branch_18_in2_data}, branch_18_in1_data}), .valid_in_bus({branch_18_in2_valid, branch_18_in1_valid}), .ready_in_bus({branch_18_in2_ready, branch_18_in1_ready}), .data_out_bus({branch_18_out2_data, branch_18_out1_data}), .valid_out_bus({branch_18_out2_valid, branch_18_out1_valid}), .ready_out_bus({branch_18_out2_ready, branch_18_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_28 (.clk(forkC_28_clk), .rst(forkC_28_rst), .data_in_bus({forkC_28_in1_data}), .valid_in_bus({forkC_28_in1_valid}), .ready_in_bus({forkC_28_in1_ready}), .data_out_bus({forkC_28_out2_data, forkC_28_out1_data}), .valid_out_bus({forkC_28_out2_valid, forkC_28_out1_valid}), .ready_out_bus({forkC_28_out2_ready, forkC_28_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) const_node_cst_3 (.clk(cst_3_clk), .rst(cst_3_rst), .data_in_bus({32'd4294967295}), .valid_in_bus({cst_3_in1_valid}), .ready_in_bus({cst_3_in1_ready}), .data_out_bus({cst_3_out1_data}), .valid_out_bus({cst_3_out1_valid}), .ready_out_bus({cst_3_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_17 (.clk(fork_17_clk), .rst(fork_17_rst), .data_in_bus({fork_17_in1_data}), .valid_in_bus({fork_17_in1_valid}), .ready_in_bus({fork_17_in1_ready}), .data_out_bus({fork_17_out5_data, fork_17_out4_data, fork_17_out3_data, fork_17_out2_data, fork_17_out1_data}), .valid_out_bus({fork_17_out5_valid, fork_17_out4_valid, fork_17_out3_valid, fork_17_out2_valid, fork_17_out1_valid}), .ready_out_bus({fork_17_out5_ready, fork_17_out4_ready, fork_17_out3_ready, fork_17_out2_ready, fork_17_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_2 (.clk(cst_2_clk), .rst(cst_2_rst), .data_in_bus({1'd0}), .valid_in_bus({cst_2_in1_valid}), .ready_in_bus({cst_2_in1_ready}), .data_out_bus({cst_2_out1_data}), .valid_out_bus({cst_2_out1_valid}), .ready_out_bus({cst_2_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block2 (.clk(brCst_block2_clk), .rst(brCst_block2_rst), .data_in_bus({1'd1}), .valid_in_bus({brCst_block2_in1_valid}), .ready_in_bus({brCst_block2_in1_ready}), .data_out_bus({brCst_block2_out1_data}), .valid_out_bus({brCst_block2_out1_valid}), .ready_out_bus({brCst_block2_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_26 (.clk(branchC_26_clk), .rst(branchC_26_rst), .data_in_bus({{branchC_26_in2_data}, branchC_26_in1_data}), .valid_in_bus({branchC_26_in2_valid, branchC_26_in1_valid}), .ready_in_bus({branchC_26_in2_ready, branchC_26_in1_ready}), .data_out_bus({branchC_26_out2_data, branchC_26_out1_data}), .valid_out_bus({branchC_26_out2_valid, branchC_26_out1_valid}), .ready_out_bus({branchC_26_out2_ready, branchC_26_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_0 (.clk(sink_0_clk), .rst(sink_0_rst), .data_in_bus({sink_0_in1_data}), .valid_in_bus({sink_0_in1_valid}), .ready_in_bus({sink_0_in1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_6 (.clk(cst_6_clk), .rst(cst_6_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_6_in1_valid}), .ready_in_bus({cst_6_in1_ready}), .data_out_bus({cst_6_out1_data}), .valid_out_bus({cst_6_out1_valid}), .ready_out_bus({cst_6_out1_ready}));
icmp_slt_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(1)) icmp_slt_op_icmp_28 (.clk(icmp_28_clk), .rst(icmp_28_rst), .data_in_bus({icmp_28_in2_data, icmp_28_in1_data}), .valid_in_bus({icmp_28_in2_valid, icmp_28_in1_valid}), .ready_in_bus({icmp_28_in2_ready, icmp_28_in1_ready}), .data_out_bus({icmp_28_out1_data}), .valid_out_bus({icmp_28_out1_valid}), .ready_out_bus({icmp_28_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) branch_node_branch_17 (.clk(branch_17_clk), .rst(branch_17_rst), .data_in_bus({{30'b0, branch_17_in2_data}, branch_17_in1_data}), .valid_in_bus({branch_17_in2_valid, branch_17_in1_valid}), .ready_in_bus({branch_17_in2_ready, branch_17_in1_ready}), .data_out_bus({branch_17_out2_data, branch_17_out1_data}), .valid_out_bus({branch_17_out2_valid, branch_17_out1_valid}), .ready_out_bus({branch_17_out2_ready, branch_17_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) branch_node_branch_19 (.clk(branch_19_clk), .rst(branch_19_rst), .data_in_bus({{30'b0, branch_19_in2_data}, branch_19_in1_data}), .valid_in_bus({branch_19_in2_valid, branch_19_in1_valid}), .ready_in_bus({branch_19_in2_ready, branch_19_in1_ready}), .data_out_bus({branch_19_out2_data, branch_19_out1_data}), .valid_out_bus({branch_19_out2_valid, branch_19_out1_valid}), .ready_out_bus({branch_19_out2_ready, branch_19_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_50 (.clk(Buffer_50_clk), .rst(Buffer_50_rst), .data_in_bus({Buffer_50_in1_data}), .valid_in_bus({Buffer_50_in1_valid}), .ready_in_bus({Buffer_50_in1_ready}), .data_out_bus({Buffer_50_out1_data}), .valid_out_bus({Buffer_50_out1_valid}), .ready_out_bus({Buffer_50_out1_ready}));
start_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) start_node_start_0 (.clk(start_0_clk), .rst(start_0_rst), .data_in_bus({start_0_in1_data}), .valid_in_bus({start_0_in1_valid}), .ready_in_bus({start_0_in1_ready}), .data_out_bus({start_0_out1_data}), .valid_out_bus({start_0_out1_valid}), .ready_out_bus({start_0_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_23 (.clk(phiC_23_clk), .rst(phiC_23_rst), .data_in_bus({phiC_23_in2_data, phiC_23_in1_data}), .valid_in_bus({phiC_23_in2_valid, phiC_23_in1_valid}), .ready_in_bus({phiC_23_in2_ready, phiC_23_in1_ready}), .data_out_bus({phiC_23_out1_data}), .valid_out_bus({phiC_23_out1_valid}), .ready_out_bus({phiC_23_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) branch_node_branch_13 (.clk(branch_13_clk), .rst(branch_13_rst), .data_in_bus({{30'b0, branch_13_in2_data}, branch_13_in1_data}), .valid_in_bus({branch_13_in2_valid, branch_13_in1_valid}), .ready_in_bus({branch_13_in2_ready, branch_13_in1_ready}), .data_out_bus({branch_13_out2_data, branch_13_out1_data}), .valid_out_bus({branch_13_out2_valid, branch_13_out1_valid}), .ready_out_bus({branch_13_out2_ready, branch_13_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) merge_node_phi_n11 (.clk(phi_n11_clk), .rst(phi_n11_rst), .data_in_bus({phi_n11_in1_data}), .valid_in_bus({phi_n11_in1_valid}), .ready_in_bus({phi_n11_in1_ready}), .data_out_bus({phi_n11_out1_data}), .valid_out_bus({phi_n11_out1_valid}), .ready_out_bus({phi_n11_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_55 (.clk(Buffer_55_clk), .rst(Buffer_55_rst), .data_in_bus({Buffer_55_in1_data}), .valid_in_bus({Buffer_55_in1_valid}), .ready_in_bus({Buffer_55_in1_ready}), .data_out_bus({Buffer_55_out1_data}), .valid_out_bus({Buffer_55_out1_valid}), .ready_out_bus({Buffer_55_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_20 (.clk(branch_20_clk), .rst(branch_20_rst), .data_in_bus({{31'b0, branch_20_in2_data}, branch_20_in1_data}), .valid_in_bus({branch_20_in2_valid, branch_20_in1_valid}), .ready_in_bus({branch_20_in2_ready, branch_20_in1_ready}), .data_out_bus({branch_20_out2_data, branch_20_out1_data}), .valid_out_bus({branch_20_out2_valid, branch_20_out1_valid}), .ready_out_bus({branch_20_out2_ready, branch_20_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n12 (.clk(phi_n12_clk), .rst(phi_n12_rst), .data_in_bus({phi_n12_in1_data}), .valid_in_bus({phi_n12_in1_valid}), .ready_in_bus({phi_n12_in1_ready}), .data_out_bus({phi_n12_out1_data}), .valid_out_bus({phi_n12_out1_valid}), .ready_out_bus({phi_n12_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_24 (.clk(forkC_24_clk), .rst(forkC_24_rst), .data_in_bus({forkC_24_in1_data}), .valid_in_bus({forkC_24_in1_valid}), .ready_in_bus({forkC_24_in1_ready}), .data_out_bus({forkC_24_out2_data, forkC_24_out1_data}), .valid_out_bus({forkC_24_out2_valid, forkC_24_out1_valid}), .ready_out_bus({forkC_24_out2_ready, forkC_24_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_12 (.clk(branch_12_clk), .rst(branch_12_rst), .data_in_bus({{31'b0, branch_12_in2_data}, branch_12_in1_data}), .valid_in_bus({branch_12_in2_valid, branch_12_in1_valid}), .ready_in_bus({branch_12_in2_ready, branch_12_in1_ready}), .data_out_bus({branch_12_out2_data, branch_12_out1_data}), .valid_out_bus({branch_12_out2_valid, branch_12_out1_valid}), .ready_out_bus({branch_12_out2_ready, branch_12_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_1 (.clk(branch_1_clk), .rst(branch_1_rst), .data_in_bus({{branch_1_in2_data}, branch_1_in1_data}), .valid_in_bus({branch_1_in2_valid, branch_1_in1_valid}), .ready_in_bus({branch_1_in2_ready, branch_1_in1_ready}), .data_out_bus({branch_1_out2_data, branch_1_out1_data}), .valid_out_bus({branch_1_out2_valid, branch_1_out1_valid}), .ready_out_bus({branch_1_out2_ready, branch_1_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_21 (.clk(phiC_21_clk), .rst(phiC_21_rst), .data_in_bus({phiC_21_in1_data}), .valid_in_bus({phiC_21_in1_valid}), .ready_in_bus({phiC_21_in1_ready}), .data_out_bus({phiC_21_out1_data}), .valid_out_bus({phiC_21_out1_valid}), .ready_out_bus({phiC_21_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_4 (.clk(branch_4_clk), .rst(branch_4_rst), .data_in_bus({{31'b0, branch_4_in2_data}, branch_4_in1_data}), .valid_in_bus({branch_4_in2_valid, branch_4_in1_valid}), .ready_in_bus({branch_4_in2_ready, branch_4_in1_ready}), .data_out_bus({branch_4_out2_data, branch_4_out1_data}), .valid_out_bus({branch_4_out2_valid, branch_4_out1_valid}), .ready_out_bus({branch_4_out2_ready, branch_4_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n14 (.clk(phi_n14_clk), .rst(phi_n14_rst), .data_in_bus({phi_n14_in1_data}), .valid_in_bus({phi_n14_in1_valid}), .ready_in_bus({phi_n14_in1_ready}), .data_out_bus({phi_n14_out1_data}), .valid_out_bus({phi_n14_out1_valid}), .ready_out_bus({phi_n14_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_10 (.clk(branch_10_clk), .rst(branch_10_rst), .data_in_bus({{31'b0, branch_10_in2_data}, branch_10_in1_data}), .valid_in_bus({branch_10_in2_valid, branch_10_in1_valid}), .ready_in_bus({branch_10_in2_ready, branch_10_in1_ready}), .data_out_bus({branch_10_out2_data, branch_10_out1_data}), .valid_out_bus({branch_10_out2_valid, branch_10_out1_valid}), .ready_out_bus({branch_10_out2_ready, branch_10_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(31))sink_node_sink_11 (.clk(sink_11_clk), .rst(sink_11_rst), .data_in_bus({sink_11_in1_data}), .valid_in_bus({sink_11_in1_valid}), .ready_in_bus({sink_11_in1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n13 (.clk(phi_n13_clk), .rst(phi_n13_rst), .data_in_bus({phi_n13_in1_data}), .valid_in_bus({phi_n13_in1_valid}), .ready_in_bus({phi_n13_in1_ready}), .data_out_bus({phi_n13_out1_data}), .valid_out_bus({phi_n13_out1_valid}), .ready_out_bus({phi_n13_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(32))source_node_source_2 (.clk(source_2_clk), .rst(source_2_rst), .data_out_bus({source_2_out1_data}), .valid_out_bus({source_2_out1_valid}), .ready_out_bus({source_2_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_7 (.clk(branch_7_clk), .rst(branch_7_rst), .data_in_bus({{31'b0, branch_7_in2_data}, branch_7_in1_data}), .valid_in_bus({branch_7_in2_valid, branch_7_in1_valid}), .ready_in_bus({branch_7_in2_ready, branch_7_in1_ready}), .data_out_bus({branch_7_out2_data, branch_7_out1_data}), .valid_out_bus({branch_7_out2_valid, branch_7_out1_valid}), .ready_out_bus({branch_7_out2_ready, branch_7_out1_ready}));
icmp_sgt_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(1)) icmp_sgt_op_icmp_9 (.clk(icmp_9_clk), .rst(icmp_9_rst), .data_in_bus({icmp_9_in2_data, icmp_9_in1_data}), .valid_in_bus({icmp_9_in2_valid, icmp_9_in1_valid}), .ready_in_bus({icmp_9_in2_ready, icmp_9_in1_ready}), .data_out_bus({icmp_9_out1_data}), .valid_out_bus({icmp_9_out1_valid}), .ready_out_bus({icmp_9_out1_ready}));
mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_8 (.clk(phi_8_clk), .rst(phi_8_rst), .data_in_bus({{31'b0, phi_8_in1_data}, phi_8_in3_data, phi_8_in2_data}), .valid_in_bus({phi_8_in1_valid, phi_8_in3_valid, phi_8_in2_valid}), .ready_in_bus({phi_8_in1_ready, phi_8_in3_ready, phi_8_in2_ready}), .data_out_bus({phi_8_out1_data}), .valid_out_bus({phi_8_out1_valid}), .ready_out_bus({phi_8_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_15 (.clk(fork_15_clk), .rst(fork_15_rst), .data_in_bus({fork_15_in1_data}), .valid_in_bus({fork_15_in1_valid}), .ready_in_bus({fork_15_in1_ready}), .data_out_bus({fork_15_out5_data, fork_15_out4_data, fork_15_out3_data, fork_15_out2_data, fork_15_out1_data}), .valid_out_bus({fork_15_out5_valid, fork_15_out4_valid, fork_15_out3_valid, fork_15_out2_valid, fork_15_out1_valid}), .ready_out_bus({fork_15_out5_ready, fork_15_out4_ready, fork_15_out3_ready, fork_15_out2_ready, fork_15_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_19 (.clk(fork_19_clk), .rst(fork_19_rst), .data_in_bus({fork_19_in1_data}), .valid_in_bus({fork_19_in1_valid}), .ready_in_bus({fork_19_in1_ready}), .data_out_bus({fork_19_out3_data, fork_19_out2_data, fork_19_out1_data}), .valid_out_bus({fork_19_out3_valid, fork_19_out2_valid, fork_19_out1_valid}), .ready_out_bus({fork_19_out3_ready, fork_19_out2_ready, fork_19_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_7 (.clk(sink_7_clk), .rst(sink_7_rst), .data_in_bus({sink_7_in1_data}), .valid_in_bus({sink_7_in1_valid}), .ready_in_bus({sink_7_in1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n9 (.clk(phi_n9_clk), .rst(phi_n9_rst), .data_in_bus({phi_n9_in1_data}), .valid_in_bus({phi_n9_in1_valid}), .ready_in_bus({phi_n9_in1_ready}), .data_out_bus({phi_n9_out1_data}), .valid_out_bus({phi_n9_out1_valid}), .ready_out_bus({phi_n9_out1_ready}));
end_node #(.INPUTS(1), .OUTPUTS(1), .MEMORY_INPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) end_node_end_0 (.clk(end_0_clk), .rst(end_0_rst), .data_in_bus({end_0_in2_data}), .valid_in_bus({end_0_in2_valid}), .ready_in_bus({end_0_in2_ready}), .e_valid_bus({end_0_in1_valid}), .e_ready_bus({end_0_in1_ready}), .data_out_bus({end_0_out1_data}), .valid_out_bus({end_0_out1_valid}), .ready_out_bus({end_0_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_15 (.clk(sink_15_clk), .rst(sink_15_rst), .data_in_bus({sink_15_in1_data}), .valid_in_bus({sink_15_in1_valid}), .ready_in_bus({sink_15_in1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) fork_node_fork_3 (.clk(fork_3_clk), .rst(fork_3_rst), .data_in_bus({fork_3_in1_data}), .valid_in_bus({fork_3_in1_valid}), .ready_in_bus({fork_3_in1_ready}), .data_out_bus({fork_3_out2_data, fork_3_out1_data}), .valid_out_bus({fork_3_out2_valid, fork_3_out1_valid}), .ready_out_bus({fork_3_out2_ready, fork_3_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_8 (.clk(fork_8_clk), .rst(fork_8_rst), .data_in_bus({fork_8_in1_data}), .valid_in_bus({fork_8_in1_valid}), .ready_in_bus({fork_8_in1_ready}), .data_out_bus({fork_8_out3_data, fork_8_out2_data, fork_8_out1_data}), .valid_out_bus({fork_8_out3_valid, fork_8_out2_valid, fork_8_out1_valid}), .ready_out_bus({fork_8_out3_ready, fork_8_out2_ready, fork_8_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_12 (.clk(sink_12_clk), .rst(sink_12_rst), .data_in_bus({sink_12_in1_data}), .valid_in_bus({sink_12_in1_valid}), .ready_in_bus({sink_12_in1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_13 (.clk(sink_13_clk), .rst(sink_13_rst), .data_in_bus({sink_13_in1_data}), .valid_in_bus({sink_13_in1_valid}), .ready_in_bus({sink_13_in1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(32))source_node_source_4 (.clk(source_4_clk), .rst(source_4_rst), .data_out_bus({source_4_out1_data}), .valid_out_bus({source_4_out1_valid}), .ready_out_bus({source_4_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_3 (.clk(branch_3_clk), .rst(branch_3_rst), .data_in_bus({{31'b0, branch_3_in2_data}, branch_3_in1_data}), .valid_in_bus({branch_3_in2_valid, branch_3_in1_valid}), .ready_in_bus({branch_3_in2_ready, branch_3_in1_ready}), .data_out_bus({branch_3_out2_data, branch_3_out1_data}), .valid_out_bus({branch_3_out2_valid, branch_3_out1_valid}), .ready_out_bus({branch_3_out2_ready, branch_3_out1_ready}));
icmp_slt_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(1)) icmp_slt_op_icmp_0 (.clk(icmp_0_clk), .rst(icmp_0_rst), .data_in_bus({icmp_0_in2_data, icmp_0_in1_data}), .valid_in_bus({icmp_0_in2_valid, icmp_0_in1_valid}), .ready_in_bus({icmp_0_in2_ready, icmp_0_in1_ready}), .data_out_bus({icmp_0_out1_data}), .valid_out_bus({icmp_0_out1_valid}), .ready_out_bus({icmp_0_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_21 (.clk(branchC_21_clk), .rst(branchC_21_rst), .data_in_bus({{branchC_21_in2_data}, branchC_21_in1_data}), .valid_in_bus({branchC_21_in2_valid, branchC_21_in1_valid}), .ready_in_bus({branchC_21_in2_ready, branchC_21_in1_ready}), .data_out_bus({branchC_21_out2_data, branchC_21_out1_data}), .valid_out_bus({branchC_21_out2_valid, branchC_21_out1_valid}), .ready_out_bus({branchC_21_out2_ready, branchC_21_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_10 (.clk(sink_10_clk), .rst(sink_10_rst), .data_in_bus({sink_10_in1_data}), .valid_in_bus({sink_10_in1_valid}), .ready_in_bus({sink_10_in1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) merge_node_phi_n7 (.clk(phi_n7_clk), .rst(phi_n7_rst), .data_in_bus({phi_n7_in2_data, phi_n7_in1_data}), .valid_in_bus({phi_n7_in2_valid, phi_n7_in1_valid}), .ready_in_bus({phi_n7_in2_ready, phi_n7_in1_ready}), .data_out_bus({phi_n7_out1_data}), .valid_out_bus({phi_n7_out1_valid}), .ready_out_bus({phi_n7_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_17 (.clk(add_17_clk), .rst(add_17_rst), .data_in_bus({add_17_in2_data, add_17_in1_data}), .valid_in_bus({add_17_in2_valid, add_17_in1_valid}), .ready_in_bus({add_17_in2_ready, add_17_in1_ready}), .data_out_bus({add_17_out1_data}), .valid_out_bus({add_17_out1_valid}), .ready_out_bus({add_17_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) OEHB_Buffer_57 (.clk(Buffer_57_clk), .rst(Buffer_57_rst), .data_in_bus({Buffer_57_in1_data}), .valid_in_bus({Buffer_57_in1_valid}), .ready_in_bus({Buffer_57_in1_ready}), .data_out_bus({Buffer_57_out1_data}), .valid_out_bus({Buffer_57_out1_valid}), .ready_out_bus({Buffer_57_out1_ready}));
icmp_sgt_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(1)) icmp_sgt_op_icmp_15 (.clk(icmp_15_clk), .rst(icmp_15_rst), .data_in_bus({icmp_15_in2_data, icmp_15_in1_data}), .valid_in_bus({icmp_15_in2_valid, icmp_15_in1_valid}), .ready_in_bus({icmp_15_in2_ready, icmp_15_in1_ready}), .data_out_bus({icmp_15_out1_data}), .valid_out_bus({icmp_15_out1_valid}), .ready_out_bus({icmp_15_out1_ready}));
start_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) start_node_n (.clk(n_clk), .rst(n_rst), .data_in_bus({n_in1_data}), .valid_in_bus({n_in1_valid}), .ready_in_bus({n_in1_ready}), .data_out_bus({n_out1_data}), .valid_out_bus({n_out1_valid}), .ready_out_bus({n_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(32), .DATA_SIZE(32)) mc_load_op_load_20 (.clk(load_20_clk), .rst(load_20_rst), .data_in_bus({load_20_in1_data}), .address_in_bus({load_20_in2_data}), .valid_in_bus({load_20_in2_valid, load_20_in1_valid}), .ready_in_bus({load_20_in2_ready, load_20_in1_ready}), .data_out_bus({load_20_out1_data}), .address_out_bus({load_20_out2_data}), .valid_out_bus({load_20_out2_valid, load_20_out1_valid}), .ready_out_bus({load_20_out2_ready, load_20_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_14 (.clk(branch_14_clk), .rst(branch_14_rst), .data_in_bus({{31'b0, branch_14_in2_data}, branch_14_in1_data}), .valid_in_bus({branch_14_in2_valid, branch_14_in1_valid}), .ready_in_bus({branch_14_in2_ready, branch_14_in1_ready}), .data_out_bus({branch_14_out2_data, branch_14_out1_data}), .valid_out_bus({branch_14_out2_valid, branch_14_out1_valid}), .ready_out_bus({branch_14_out2_ready, branch_14_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_14 (.clk(sink_14_clk), .rst(sink_14_rst), .data_in_bus({sink_14_in1_data}), .valid_in_bus({sink_14_in1_valid}), .ready_in_bus({sink_14_in1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) const_node_cst_4 (.clk(cst_4_clk), .rst(cst_4_rst), .data_in_bus({32'd4294967295}), .valid_in_bus({cst_4_in1_valid}), .ready_in_bus({cst_4_in1_ready}), .data_out_bus({cst_4_out1_data}), .valid_out_bus({cst_4_out1_valid}), .ready_out_bus({cst_4_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(32))source_node_source_3 (.clk(source_3_clk), .rst(source_3_rst), .data_out_bus({source_3_out1_data}), .valid_out_bus({source_3_out1_valid}), .ready_out_bus({source_3_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) branch_node_branch_5 (.clk(branch_5_clk), .rst(branch_5_rst), .data_in_bus({{30'b0, branch_5_in2_data}, branch_5_in1_data}), .valid_in_bus({branch_5_in2_valid, branch_5_in1_valid}), .ready_in_bus({branch_5_in2_ready, branch_5_in1_ready}), .data_out_bus({branch_5_out2_data, branch_5_out1_data}), .valid_out_bus({branch_5_out2_valid, branch_5_out1_valid}), .ready_out_bus({branch_5_out2_ready, branch_5_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_1 (.clk(sink_1_clk), .rst(sink_1_rst), .data_in_bus({sink_1_in1_data}), .valid_in_bus({sink_1_in1_valid}), .ready_in_bus({sink_1_in1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_27 (.clk(branchC_27_clk), .rst(branchC_27_rst), .data_in_bus({{branchC_27_in2_data}, branchC_27_in1_data}), .valid_in_bus({branchC_27_in2_valid, branchC_27_in1_valid}), .ready_in_bus({branchC_27_in2_ready, branchC_27_in1_ready}), .data_out_bus({branchC_27_out2_data, branchC_27_out1_data}), .valid_out_bus({branchC_27_out2_valid, branchC_27_out1_valid}), .ready_out_bus({branchC_27_out2_ready, branchC_27_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_2 (.clk(sink_2_clk), .rst(sink_2_rst), .data_in_bus({sink_2_in1_data}), .valid_in_bus({sink_2_in1_valid}), .ready_in_bus({sink_2_in1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_25 (.clk(branchC_25_clk), .rst(branchC_25_rst), .data_in_bus({{branchC_25_in2_data}, branchC_25_in1_data}), .valid_in_bus({branchC_25_in2_valid, branchC_25_in1_valid}), .ready_in_bus({branchC_25_in2_ready, branchC_25_in1_ready}), .data_out_bus({branchC_25_out2_data, branchC_25_out1_data}), .valid_out_bus({branchC_25_out2_valid, branchC_25_out1_valid}), .ready_out_bus({branchC_25_out2_ready, branchC_25_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_4 (.clk(fork_4_clk), .rst(fork_4_rst), .data_in_bus({fork_4_in1_data}), .valid_in_bus({fork_4_in1_valid}), .ready_in_bus({fork_4_in1_ready}), .data_out_bus({fork_4_out2_data, fork_4_out1_data}), .valid_out_bus({fork_4_out2_valid, fork_4_out1_valid}), .ready_out_bus({fork_4_out2_ready, fork_4_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_22 (.clk(fork_22_clk), .rst(fork_22_rst), .data_in_bus({fork_22_in1_data}), .valid_in_bus({fork_22_in1_valid}), .ready_in_bus({fork_22_in1_ready}), .data_out_bus({fork_22_out2_data, fork_22_out1_data}), .valid_out_bus({fork_22_out2_valid, fork_22_out1_valid}), .ready_out_bus({fork_22_out2_ready, fork_22_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_51 (.clk(Buffer_51_clk), .rst(Buffer_51_rst), .data_in_bus({Buffer_51_in1_data}), .valid_in_bus({Buffer_51_in1_valid}), .ready_in_bus({Buffer_51_in1_ready}), .data_out_bus({Buffer_51_out1_data}), .valid_out_bus({Buffer_51_out1_valid}), .ready_out_bus({Buffer_51_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n0 (.clk(phi_n0_clk), .rst(phi_n0_rst), .data_in_bus({phi_n0_in1_data}), .valid_in_bus({phi_n0_in1_valid}), .ready_in_bus({phi_n0_in1_ready}), .data_out_bus({phi_n0_out1_data}), .valid_out_bus({phi_n0_out1_valid}), .ready_out_bus({phi_n0_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_22 (.clk(phiC_22_clk), .rst(phiC_22_rst), .data_in_bus({phiC_22_in2_data, phiC_22_in1_data}), .valid_in_bus({phiC_22_in2_valid, phiC_22_in1_valid}), .ready_in_bus({phiC_22_in2_ready, phiC_22_in1_ready}), .data_out_bus({phiC_22_out1_data}), .valid_out_bus({phiC_22_out1_valid}), .ready_out_bus({phiC_22_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n1 (.clk(phi_n1_clk), .rst(phi_n1_rst), .data_in_bus({phi_n1_in2_data, phi_n1_in1_data}), .valid_in_bus({phi_n1_in2_valid, phi_n1_in1_valid}), .ready_in_bus({phi_n1_in2_ready, phi_n1_in1_ready}), .data_out_bus({phi_n1_out1_data}), .valid_out_bus({phi_n1_out1_valid}), .ready_out_bus({phi_n1_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_2 (.clk(fork_2_clk), .rst(fork_2_rst), .data_in_bus({fork_2_in1_data}), .valid_in_bus({fork_2_in1_valid}), .ready_in_bus({fork_2_in1_ready}), .data_out_bus({fork_2_out2_data, fork_2_out1_data}), .valid_out_bus({fork_2_out2_valid, fork_2_out1_valid}), .ready_out_bus({fork_2_out2_ready, fork_2_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_16 (.clk(branch_16_clk), .rst(branch_16_rst), .data_in_bus({{31'b0, branch_16_in2_data}, branch_16_in1_data}), .valid_in_bus({branch_16_in2_valid, branch_16_in1_valid}), .ready_in_bus({branch_16_in2_ready, branch_16_in1_ready}), .data_out_bus({branch_16_out2_data, branch_16_out1_data}), .valid_out_bus({branch_16_out2_valid, branch_16_out1_valid}), .ready_out_bus({branch_16_out2_ready, branch_16_out1_ready}));
ret_op #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) ret_op_ret_0 (.clk(ret_0_clk), .rst(ret_0_rst), .data_in_bus({ret_0_in1_data}), .valid_in_bus({ret_0_in1_valid}), .ready_in_bus({ret_0_in1_ready}), .data_out_bus({ret_0_out1_data}), .valid_out_bus({ret_0_out1_valid}), .ready_out_bus({ret_0_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) OEHB_Buffer_52 (.clk(Buffer_52_clk), .rst(Buffer_52_rst), .data_in_bus({Buffer_52_in1_data}), .valid_in_bus({Buffer_52_in1_valid}), .ready_in_bus({Buffer_52_in1_ready}), .data_out_bus({Buffer_52_out1_data}), .valid_out_bus({Buffer_52_out1_valid}), .ready_out_bus({Buffer_52_out1_ready}));
mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31), .COND_SIZE(1)) mux_node_phi_3 (.clk(phi_3_clk), .rst(phi_3_rst), .data_in_bus({{30'b0, phi_3_in1_data}, phi_3_in3_data, phi_3_in2_data}), .valid_in_bus({phi_3_in1_valid, phi_3_in3_valid, phi_3_in2_valid}), .ready_in_bus({phi_3_in1_ready, phi_3_in3_ready, phi_3_in2_ready}), .data_out_bus({phi_3_out1_data}), .valid_out_bus({phi_3_out1_valid}), .ready_out_bus({phi_3_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_8 (.clk(branch_8_clk), .rst(branch_8_rst), .data_in_bus({{31'b0, branch_8_in2_data}, branch_8_in1_data}), .valid_in_bus({branch_8_in2_valid, branch_8_in1_valid}), .ready_in_bus({branch_8_in2_ready, branch_8_in1_ready}), .data_out_bus({branch_8_out2_data, branch_8_out1_data}), .valid_out_bus({branch_8_out2_valid, branch_8_out1_valid}), .ready_out_bus({branch_8_out2_ready, branch_8_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_5 (.clk(source_5_clk), .rst(source_5_rst), .data_out_bus({source_5_out1_data}), .valid_out_bus({source_5_out1_valid}), .ready_out_bus({source_5_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_8 (.clk(sink_8_clk), .rst(sink_8_rst), .data_in_bus({sink_8_in1_data}), .valid_in_bus({sink_8_in1_valid}), .ready_in_bus({sink_8_in1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_3 (.clk(sink_3_clk), .rst(sink_3_rst), .data_in_bus({sink_3_in1_data}), .valid_in_bus({sink_3_in1_valid}), .ready_in_bus({sink_3_in1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_53 (.clk(Buffer_53_clk), .rst(Buffer_53_rst), .data_in_bus({Buffer_53_in1_data}), .valid_in_bus({Buffer_53_in1_valid}), .ready_in_bus({Buffer_53_in1_ready}), .data_out_bus({Buffer_53_out1_data}), .valid_out_bus({Buffer_53_out1_valid}), .ready_out_bus({Buffer_53_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n16 (.clk(phi_n16_clk), .rst(phi_n16_rst), .data_in_bus({phi_n16_in1_data}), .valid_in_bus({phi_n16_in1_valid}), .ready_in_bus({phi_n16_in1_ready}), .data_out_bus({phi_n16_out1_data}), .valid_out_bus({phi_n16_out1_valid}), .ready_out_bus({phi_n16_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_11 (.clk(add_11_clk), .rst(add_11_rst), .data_in_bus({add_11_in2_data, add_11_in1_data}), .valid_in_bus({add_11_in2_valid, add_11_in1_valid}), .ready_in_bus({add_11_in2_ready, add_11_in1_ready}), .data_out_bus({add_11_out1_data}), .valid_out_bus({add_11_out1_valid}), .ready_out_bus({add_11_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_0 (.clk(fork_0_clk), .rst(fork_0_rst), .data_in_bus({fork_0_in1_data}), .valid_in_bus({fork_0_in1_valid}), .ready_in_bus({fork_0_in1_ready}), .data_out_bus({fork_0_out2_data, fork_0_out1_data}), .valid_out_bus({fork_0_out2_valid, fork_0_out1_valid}), .ready_out_bus({fork_0_out2_ready, fork_0_out1_ready}));
mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(32), .DATA_SIZE(32)) mc_store_op_store_0 (.clk(store_0_clk), .rst(store_0_rst), .data_in_bus({store_0_in1_data}), .address_in_bus({store_0_in2_data}), .valid_in_bus({store_0_in2_valid, store_0_in1_valid}), .ready_in_bus({store_0_in2_ready, store_0_in1_ready}), .data_out_bus({store_0_out1_data}), .address_out_bus({store_0_out2_data}), .valid_out_bus({store_0_out2_valid, store_0_out1_valid}), .ready_out_bus({store_0_out2_ready, store_0_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) add_op_add_27 (.clk(add_27_clk), .rst(add_27_rst), .data_in_bus({add_27_in2_data, add_27_in1_data}), .valid_in_bus({add_27_in2_valid, add_27_in1_valid}), .ready_in_bus({add_27_in2_ready, add_27_in1_ready}), .data_out_bus({add_27_out1_data}), .valid_out_bus({add_27_out1_valid}), .ready_out_bus({add_27_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_8 (.clk(cst_8_clk), .rst(cst_8_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_8_in1_valid}), .ready_in_bus({cst_8_in1_ready}), .data_out_bus({cst_8_out1_data}), .valid_out_bus({cst_8_out1_valid}), .ready_out_bus({cst_8_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(31), .DATA_SIZE(32)) mc_load_op_load_6 (.clk(load_6_clk), .rst(load_6_rst), .data_in_bus({load_6_in1_data}), .address_in_bus({load_6_in2_data}), .valid_in_bus({load_6_in2_valid, load_6_in1_valid}), .ready_in_bus({load_6_in2_ready, load_6_in1_ready}), .data_out_bus({load_6_out1_data}), .address_out_bus({load_6_out2_data}), .valid_out_bus({load_6_out2_valid, load_6_out1_valid}), .ready_out_bus({load_6_out2_ready, load_6_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_14 (.clk(fork_14_clk), .rst(fork_14_rst), .data_in_bus({fork_14_in1_data}), .valid_in_bus({fork_14_in1_valid}), .ready_in_bus({fork_14_in1_ready}), .data_out_bus({fork_14_out3_data, fork_14_out2_data, fork_14_out1_data}), .valid_out_bus({fork_14_out3_valid, fork_14_out2_valid, fork_14_out1_valid}), .ready_out_bus({fork_14_out3_ready, fork_14_out2_ready, fork_14_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block6 (.clk(brCst_block6_clk), .rst(brCst_block6_rst), .data_in_bus({1'd1}), .valid_in_bus({brCst_block6_in1_valid}), .ready_in_bus({brCst_block6_in1_ready}), .data_out_bus({brCst_block6_out1_data}), .valid_out_bus({brCst_block6_out1_valid}), .ready_out_bus({brCst_block6_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) merge_node_phi_n15 (.clk(phi_n15_clk), .rst(phi_n15_rst), .data_in_bus({phi_n15_in1_data}), .valid_in_bus({phi_n15_in1_valid}), .ready_in_bus({phi_n15_in1_ready}), .data_out_bus({phi_n15_out1_data}), .valid_out_bus({phi_n15_out1_valid}), .ready_out_bus({phi_n15_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) fork_node_fork_1 (.clk(fork_1_clk), .rst(fork_1_rst), .data_in_bus({fork_1_in1_data}), .valid_in_bus({fork_1_in1_valid}), .ready_in_bus({fork_1_in1_ready}), .data_out_bus({fork_1_out3_data, fork_1_out2_data, fork_1_out1_data}), .valid_out_bus({fork_1_out3_valid, fork_1_out2_valid, fork_1_out1_valid}), .ready_out_bus({fork_1_out3_ready, fork_1_out2_ready, fork_1_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block3 (.clk(brCst_block3_clk), .rst(brCst_block3_rst), .data_in_bus({1'd1}), .valid_in_bus({brCst_block3_in1_valid}), .ready_in_bus({brCst_block3_in1_ready}), .data_out_bus({brCst_block3_out1_data}), .valid_out_bus({brCst_block3_out1_valid}), .ready_out_bus({brCst_block3_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_20 (.clk(phiC_20_clk), .rst(phiC_20_rst), .data_in_bus({phiC_20_in1_data}), .valid_in_bus({phiC_20_in1_valid}), .ready_in_bus({phiC_20_in1_ready}), .data_out_bus({phiC_20_out1_data}), .valid_out_bus({phiC_20_out1_valid}), .ready_out_bus({phiC_20_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_0 (.clk(cst_0_clk), .rst(cst_0_rst), .data_in_bus({2'd2}), .valid_in_bus({cst_0_in1_valid}), .ready_in_bus({cst_0_in1_ready}), .data_out_bus({cst_0_out1_data}), .valid_out_bus({cst_0_out1_valid}), .ready_out_bus({cst_0_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_18 (.clk(fork_18_clk), .rst(fork_18_rst), .data_in_bus({fork_18_in1_data}), .valid_in_bus({fork_18_in1_valid}), .ready_in_bus({fork_18_in1_ready}), .data_out_bus({fork_18_out5_data, fork_18_out4_data, fork_18_out3_data, fork_18_out2_data, fork_18_out1_data}), .valid_out_bus({fork_18_out5_valid, fork_18_out4_valid, fork_18_out3_valid, fork_18_out2_valid, fork_18_out1_valid}), .ready_out_bus({fork_18_out5_ready, fork_18_out4_ready, fork_18_out3_ready, fork_18_out2_ready, fork_18_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) OEHB_Buffer_58 (.clk(Buffer_58_clk), .rst(Buffer_58_rst), .data_in_bus({Buffer_58_in1_data}), .valid_in_bus({Buffer_58_in1_valid}), .ready_in_bus({Buffer_58_in1_ready}), .data_out_bus({Buffer_58_out1_data}), .valid_out_bus({Buffer_58_out1_valid}), .ready_out_bus({Buffer_58_out1_ready}));
mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(32), .DATA_SIZE(32)) mc_store_op_store_1 (.clk(store_1_clk), .rst(store_1_rst), .data_in_bus({store_1_in1_data}), .address_in_bus({store_1_in2_data}), .valid_in_bus({store_1_in2_valid, store_1_in1_valid}), .ready_in_bus({store_1_in2_ready, store_1_in1_ready}), .data_out_bus({store_1_out1_data}), .address_out_bus({store_1_out2_data}), .valid_out_bus({store_1_out2_valid, store_1_out1_valid}), .ready_out_bus({store_1_out2_ready, store_1_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n8 (.clk(phi_n8_clk), .rst(phi_n8_rst), .data_in_bus({phi_n8_in2_data, phi_n8_in1_data}), .valid_in_bus({phi_n8_in2_valid, phi_n8_in1_valid}), .ready_in_bus({phi_n8_in2_ready, phi_n8_in1_ready}), .data_out_bus({phi_n8_out1_data}), .valid_out_bus({phi_n8_out1_valid}), .ready_out_bus({phi_n8_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_23 (.clk(forkC_23_clk), .rst(forkC_23_rst), .data_in_bus({forkC_23_in1_data}), .valid_in_bus({forkC_23_in1_valid}), .ready_in_bus({forkC_23_in1_ready}), .data_out_bus({forkC_23_out3_data, forkC_23_out2_data, forkC_23_out1_data}), .valid_out_bus({forkC_23_out3_valid, forkC_23_out2_valid, forkC_23_out1_valid}), .ready_out_bus({forkC_23_out3_ready, forkC_23_out2_ready, forkC_23_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) branch_node_branch_9 (.clk(branch_9_clk), .rst(branch_9_rst), .data_in_bus({{30'b0, branch_9_in2_data}, branch_9_in1_data}), .valid_in_bus({branch_9_in2_valid, branch_9_in1_valid}), .ready_in_bus({branch_9_in2_ready, branch_9_in1_ready}), .data_out_bus({branch_9_out2_data, branch_9_out1_data}), .valid_out_bus({branch_9_out2_valid, branch_9_out1_valid}), .ready_out_bus({branch_9_out2_ready, branch_9_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_1 (.clk(source_1_clk), .rst(source_1_rst), .data_out_bus({source_1_out1_data}), .valid_out_bus({source_1_out1_valid}), .ready_out_bus({source_1_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n5 (.clk(phi_n5_clk), .rst(phi_n5_rst), .data_in_bus({phi_n5_in2_data, phi_n5_in1_data}), .valid_in_bus({phi_n5_in2_valid, phi_n5_in1_valid}), .ready_in_bus({phi_n5_in2_ready, phi_n5_in1_ready}), .data_out_bus({phi_n5_out1_data}), .valid_out_bus({phi_n5_out1_valid}), .ready_out_bus({phi_n5_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_1 (.clk(cst_1_clk), .rst(cst_1_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_1_in1_valid}), .ready_in_bus({cst_1_in1_ready}), .data_out_bus({cst_1_out1_data}), .valid_out_bus({cst_1_out1_valid}), .ready_out_bus({cst_1_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_16 (.clk(fork_16_clk), .rst(fork_16_rst), .data_in_bus({fork_16_in1_data}), .valid_in_bus({fork_16_in1_valid}), .ready_in_bus({fork_16_in1_ready}), .data_out_bus({fork_16_out5_data, fork_16_out4_data, fork_16_out3_data, fork_16_out2_data, fork_16_out1_data}), .valid_out_bus({fork_16_out5_valid, fork_16_out4_valid, fork_16_out3_valid, fork_16_out2_valid, fork_16_out1_valid}), .ready_out_bus({fork_16_out5_ready, fork_16_out4_ready, fork_16_out3_ready, fork_16_out2_ready, fork_16_out1_ready}));
source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_0 (.clk(source_0_clk), .rst(source_0_rst), .data_out_bus({source_0_out1_data}), .valid_out_bus({source_0_out1_valid}), .ready_out_bus({source_0_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) merge_node_phi_n4 (.clk(phi_n4_clk), .rst(phi_n4_rst), .data_in_bus({phi_n4_in2_data, phi_n4_in1_data}), .valid_in_bus({phi_n4_in2_valid, phi_n4_in1_valid}), .ready_in_bus({phi_n4_in2_ready, phi_n4_in1_ready}), .data_out_bus({phi_n4_out1_data}), .valid_out_bus({phi_n4_out1_valid}), .ready_out_bus({phi_n4_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_15 (.clk(branch_15_clk), .rst(branch_15_rst), .data_in_bus({{31'b0, branch_15_in2_data}, branch_15_in1_data}), .valid_in_bus({branch_15_in2_valid, branch_15_in1_valid}), .ready_in_bus({branch_15_in2_ready, branch_15_in1_ready}), .data_out_bus({branch_15_out2_data, branch_15_out1_data}), .valid_out_bus({branch_15_out2_valid, branch_15_out1_valid}), .ready_out_bus({branch_15_out2_ready, branch_15_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_22 (.clk(branchC_22_clk), .rst(branchC_22_rst), .data_in_bus({{branchC_22_in2_data}, branchC_22_in1_data}), .valid_in_bus({branchC_22_in2_valid, branchC_22_in1_valid}), .ready_in_bus({branchC_22_in2_ready, branchC_22_in1_ready}), .data_out_bus({branchC_22_out2_data, branchC_22_out1_data}), .valid_out_bus({branchC_22_out2_valid, branchC_22_out1_valid}), .ready_out_bus({branchC_22_out2_ready, branchC_22_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_0 (.clk(branch_0_clk), .rst(branch_0_rst), .data_in_bus({{31'b0, branch_0_in2_data}, branch_0_in1_data}), .valid_in_bus({branch_0_in2_valid, branch_0_in1_valid}), .ready_in_bus({branch_0_in2_ready, branch_0_in1_ready}), .data_out_bus({branch_0_out2_data, branch_0_out1_data}), .valid_out_bus({branch_0_out2_valid, branch_0_out1_valid}), .ready_out_bus({branch_0_out2_ready, branch_0_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(31))sink_node_sink_6 (.clk(sink_6_clk), .rst(sink_6_rst), .data_in_bus({sink_6_in1_data}), .valid_in_bus({sink_6_in1_valid}), .ready_in_bus({sink_6_in1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_23 (.clk(branchC_23_clk), .rst(branchC_23_rst), .data_in_bus({{branchC_23_in2_data}, branchC_23_in1_data}), .valid_in_bus({branchC_23_in2_valid, branchC_23_in1_valid}), .ready_in_bus({branchC_23_in2_ready, branchC_23_in1_ready}), .data_out_bus({branchC_23_out2_data, branchC_23_out1_data}), .valid_out_bus({branchC_23_out2_valid, branchC_23_out1_valid}), .ready_out_bus({branchC_23_out2_ready, branchC_23_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_11 (.clk(branch_11_clk), .rst(branch_11_rst), .data_in_bus({{31'b0, branch_11_in2_data}, branch_11_in1_data}), .valid_in_bus({branch_11_in2_valid, branch_11_in1_valid}), .ready_in_bus({branch_11_in2_ready, branch_11_in1_ready}), .data_out_bus({branch_11_out2_data, branch_11_out1_data}), .valid_out_bus({branch_11_out2_valid, branch_11_out1_valid}), .ready_out_bus({branch_11_out2_ready, branch_11_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n2 (.clk(phi_n2_clk), .rst(phi_n2_rst), .data_in_bus({phi_n2_in2_data, phi_n2_in1_data}), .valid_in_bus({phi_n2_in2_valid, phi_n2_in1_valid}), .ready_in_bus({phi_n2_in2_ready, phi_n2_in1_ready}), .data_out_bus({phi_n2_out1_data}), .valid_out_bus({phi_n2_out1_valid}), .ready_out_bus({phi_n2_out1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) OEHB_Buffer_56 (.clk(Buffer_56_clk), .rst(Buffer_56_rst), .data_in_bus({Buffer_56_in1_data}), .valid_in_bus({Buffer_56_in1_valid}), .ready_in_bus({Buffer_56_in1_ready}), .data_out_bus({Buffer_56_out1_data}), .valid_out_bus({Buffer_56_out1_valid}), .ready_out_bus({Buffer_56_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_27 (.clk(forkC_27_clk), .rst(forkC_27_rst), .data_in_bus({forkC_27_in1_data}), .valid_in_bus({forkC_27_in1_valid}), .ready_in_bus({forkC_27_in1_ready}), .data_out_bus({forkC_27_out3_data, forkC_27_out2_data, forkC_27_out1_data}), .valid_out_bus({forkC_27_out3_valid, forkC_27_out2_valid, forkC_27_out1_valid}), .ready_out_bus({forkC_27_out3_ready, forkC_27_out2_ready, forkC_27_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n3 (.clk(phi_n3_clk), .rst(phi_n3_rst), .data_in_bus({phi_n3_in2_data, phi_n3_in1_data}), .valid_in_bus({phi_n3_in2_valid, phi_n3_in1_valid}), .ready_in_bus({phi_n3_in2_ready, phi_n3_in1_ready}), .data_out_bus({phi_n3_out1_data}), .valid_out_bus({phi_n3_out1_valid}), .ready_out_bus({phi_n3_out1_ready}));
add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_23 (.clk(add_23_clk), .rst(add_23_rst), .data_in_bus({add_23_in2_data, add_23_in1_data}), .valid_in_bus({add_23_in2_valid, add_23_in1_valid}), .ready_in_bus({add_23_in2_ready, add_23_in1_ready}), .data_out_bus({add_23_out1_data}), .valid_out_bus({add_23_out1_valid}), .ready_out_bus({add_23_out1_ready}));
cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_18 (.clk(phiC_18_clk), .rst(phiC_18_rst), .data_in_bus({phiC_18_in2_data, phiC_18_in1_data}), .valid_in_bus({phiC_18_in2_valid, phiC_18_in1_valid}), .ready_in_bus({phiC_18_in2_ready, phiC_18_in1_ready}), .data_out_bus({phiC_18_out2_data, phiC_18_out1_data}), .valid_out_bus({phiC_18_out2_valid, phiC_18_out1_valid}), .ready_out_bus({phiC_18_out2_ready, phiC_18_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_7 (.clk(cst_7_clk), .rst(cst_7_rst), .data_in_bus({1'd1}), .valid_in_bus({cst_7_in1_valid}), .ready_in_bus({cst_7_in1_ready}), .data_out_bus({cst_7_out1_data}), .valid_out_bus({cst_7_out1_valid}), .ready_out_bus({cst_7_out1_ready}));
const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) const_node_cst_5 (.clk(cst_5_clk), .rst(cst_5_rst), .data_in_bus({32'd4294967295}), .valid_in_bus({cst_5_in1_valid}), .ready_in_bus({cst_5_in1_ready}), .data_out_bus({cst_5_out1_data}), .valid_out_bus({cst_5_out1_valid}), .ready_out_bus({cst_5_out1_ready}));
merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n6 (.clk(phi_n6_clk), .rst(phi_n6_rst), .data_in_bus({phi_n6_in2_data, phi_n6_in1_data}), .valid_in_bus({phi_n6_in2_valid, phi_n6_in1_valid}), .ready_in_bus({phi_n6_in2_ready, phi_n6_in1_ready}), .data_out_bus({phi_n6_out1_data}), .valid_out_bus({phi_n6_out1_valid}), .ready_out_bus({phi_n6_out1_ready}));
mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(32), .DATA_SIZE(32)) mc_load_op_load_14 (.clk(load_14_clk), .rst(load_14_rst), .data_in_bus({load_14_in1_data}), .address_in_bus({load_14_in2_data}), .valid_in_bus({load_14_in2_valid, load_14_in1_valid}), .ready_in_bus({load_14_in2_ready, load_14_in1_ready}), .data_out_bus({load_14_out1_data}), .address_out_bus({load_14_out2_data}), .valid_out_bus({load_14_out2_valid, load_14_out1_valid}), .ready_out_bus({load_14_out2_ready, load_14_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(31))sink_node_sink_9 (.clk(sink_9_clk), .rst(sink_9_rst), .data_in_bus({sink_9_in1_data}), .valid_in_bus({sink_9_in1_valid}), .ready_in_bus({sink_9_in1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) branch_node_branch_6 (.clk(branch_6_clk), .rst(branch_6_rst), .data_in_bus({{30'b0, branch_6_in2_data}, branch_6_in1_data}), .valid_in_bus({branch_6_in2_valid, branch_6_in1_valid}), .ready_in_bus({branch_6_in2_ready, branch_6_in1_ready}), .data_out_bus({branch_6_out2_data, branch_6_out1_data}), .valid_out_bus({branch_6_out2_valid, branch_6_out1_valid}), .ready_out_bus({branch_6_out2_ready, branch_6_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_4 (.clk(sink_4_clk), .rst(sink_4_rst), .data_in_bus({sink_4_in1_data}), .valid_in_bus({sink_4_in1_valid}), .ready_in_bus({sink_4_in1_ready}));
OEHB #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(31), .DATA_OUT_SIZE(31)) OEHB_Buffer_54 (.clk(Buffer_54_clk), .rst(Buffer_54_rst), .data_in_bus({Buffer_54_in1_data}), .valid_in_bus({Buffer_54_in1_valid}), .ready_in_bus({Buffer_54_in1_ready}), .data_out_bus({Buffer_54_out1_data}), .valid_out_bus({Buffer_54_out1_valid}), .ready_out_bus({Buffer_54_out1_ready}));
cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_19 (.clk(phiC_19_clk), .rst(phiC_19_rst), .data_in_bus({phiC_19_in2_data, phiC_19_in1_data}), .valid_in_bus({phiC_19_in2_valid, phiC_19_in1_valid}), .ready_in_bus({phiC_19_in2_ready, phiC_19_in1_ready}), .data_out_bus({phiC_19_out2_data, phiC_19_out1_data}), .valid_out_bus({phiC_19_out2_valid, phiC_19_out1_valid}), .ready_out_bus({phiC_19_out2_ready, phiC_19_out1_ready}));
merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n10 (.clk(phi_n10_clk), .rst(phi_n10_rst), .data_in_bus({phi_n10_in1_data}), .valid_in_bus({phi_n10_in1_valid}), .ready_in_bus({phi_n10_in1_ready}), .data_out_bus({phi_n10_out1_data}), .valid_out_bus({phi_n10_out1_valid}), .ready_out_bus({phi_n10_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_2 (.clk(branch_2_clk), .rst(branch_2_rst), .data_in_bus({{31'b0, branch_2_in2_data}, branch_2_in1_data}), .valid_in_bus({branch_2_in2_valid, branch_2_in1_valid}), .ready_in_bus({branch_2_in2_ready, branch_2_in1_ready}), .data_out_bus({branch_2_out2_data, branch_2_out1_data}), .valid_out_bus({branch_2_out2_valid, branch_2_out1_valid}), .ready_out_bus({branch_2_out2_ready, branch_2_out1_ready}));
branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_24 (.clk(branchC_24_clk), .rst(branchC_24_rst), .data_in_bus({{branchC_24_in2_data}, branchC_24_in1_data}), .valid_in_bus({branchC_24_in2_valid, branchC_24_in1_valid}), .ready_in_bus({branchC_24_in2_ready, branchC_24_in1_ready}), .data_out_bus({branchC_24_out2_data, branchC_24_out1_data}), .valid_out_bus({branchC_24_out2_valid, branchC_24_out1_valid}), .ready_out_bus({branchC_24_out2_ready, branchC_24_out1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_10 (.clk(fork_10_clk), .rst(fork_10_rst), .data_in_bus({fork_10_in1_data}), .valid_in_bus({fork_10_in1_valid}), .ready_in_bus({fork_10_in1_ready}), .data_out_bus({fork_10_out2_data, fork_10_out1_data}), .valid_out_bus({fork_10_out2_valid, fork_10_out1_valid}), .ready_out_bus({fork_10_out2_ready, fork_10_out1_ready}));
sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(31))sink_node_sink_5 (.clk(sink_5_clk), .rst(sink_5_rst), .data_in_bus({sink_5_in1_data}), .valid_in_bus({sink_5_in1_valid}), .ready_in_bus({sink_5_in1_ready}));
fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_9 (.clk(fork_9_clk), .rst(fork_9_rst), .data_in_bus({fork_9_in1_data}), .valid_in_bus({fork_9_in1_valid}), .ready_in_bus({fork_9_in1_ready}), .data_out_bus({fork_9_out2_data, fork_9_out1_data}), .valid_out_bus({fork_9_out2_valid, fork_9_out1_valid}), .ready_out_bus({fork_9_out2_ready, fork_9_out1_ready}));
endmodule
