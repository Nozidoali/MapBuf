module stencil_2d(
	input clk,
	input rst,

	output [31 : 0]end_out,
	output end_valid,
	input end_ready,

	input [0 : 0]start_in,
	input start_valid,
	output start_ready,

	output [5 : 0]filter_address0,
	output filter_ce0,
	output filter_we0,
	output [31 : 0]filter_dout0,
	input [31 : 0]filter_din0,
	output [5 : 0]filter_address1,
	output filter_ce1,
	output filter_we1,
	output [31 : 0]filter_dout1,
	input [31 : 0]filter_din1,

	output [12 : 0]orig_address0,
	output orig_ce0,
	output orig_we0,
	output [31 : 0]orig_dout0,
	input [31 : 0]orig_din0,
	output [12 : 0]orig_address1,
	output orig_ce1,
	output orig_we1,
	output [31 : 0]orig_dout1,
	input [31 : 0]orig_din1,

	output [10 : 0]sol_address0,
	output sol_ce0,
	output sol_we0,
	output [31 : 0]sol_dout0,
	input [31 : 0]sol_din0,
	output [10 : 0]sol_address1,
	output sol_ce1,
	output sol_we1,
	output [31 : 0]sol_dout1,
	input [31 : 0]sol_din1

);

	wire phi_5_clk;
	wire phi_5_rst;
	wire [0 : 0]phi_5_in1_data;
	wire phi_5_in1_ready;
	wire phi_5_in1_valid;
	wire [2 : 0]phi_5_in2_data;
	wire phi_5_in2_ready;
	wire phi_5_in2_valid;
	wire [2 : 0]phi_5_in3_data;
	wire phi_5_in3_ready;
	wire phi_5_in3_valid;
	wire [2 : 0]phi_5_out1_data;
	wire phi_5_out1_ready;
	wire phi_5_out1_valid;

	wire phi_6_clk;
	wire phi_6_rst;
	wire [0 : 0]phi_6_in1_data;
	wire phi_6_in1_ready;
	wire phi_6_in1_valid;
	wire [31 : 0]phi_6_in2_data;
	wire phi_6_in2_ready;
	wire phi_6_in2_valid;
	wire [31 : 0]phi_6_in3_data;
	wire phi_6_in3_ready;
	wire phi_6_in3_valid;
	wire [31 : 0]phi_6_out1_data;
	wire phi_6_out1_ready;
	wire phi_6_out1_valid;

	wire brCst_block4_clk;
	wire brCst_block4_rst;
	wire [0 : 0]brCst_block4_in1_data;
	wire brCst_block4_in1_ready;
	wire brCst_block4_in1_valid;
	wire [0 : 0]brCst_block4_out1_data;
	wire brCst_block4_out1_ready;
	wire brCst_block4_out1_valid;

	wire cst_4_clk;
	wire cst_4_rst;
	wire [0 : 0]cst_4_in1_data;
	wire cst_4_in1_ready;
	wire cst_4_in1_valid;
	wire [0 : 0]cst_4_out1_data;
	wire cst_4_out1_ready;
	wire cst_4_out1_valid;

	wire phi_n6_clk;
	wire phi_n6_rst;
	wire [4 : 0]phi_n6_in1_data;
	wire phi_n6_in1_ready;
	wire phi_n6_in1_valid;
	wire [4 : 0]phi_n6_in2_data;
	wire phi_n6_in2_ready;
	wire phi_n6_in2_valid;
	wire [4 : 0]phi_n6_out1_data;
	wire phi_n6_out1_ready;
	wire phi_n6_out1_valid;

	wire phi_n7_clk;
	wire phi_n7_rst;
	wire [4 : 0]phi_n7_in1_data;
	wire phi_n7_in1_ready;
	wire phi_n7_in1_valid;
	wire [4 : 0]phi_n7_in2_data;
	wire phi_n7_in2_ready;
	wire phi_n7_in2_valid;
	wire [4 : 0]phi_n7_out1_data;
	wire phi_n7_out1_ready;
	wire phi_n7_out1_valid;

	wire branch_7_clk;
	wire branch_7_rst;
	wire [0 : 0]branch_7_in1_data;
	wire branch_7_in1_ready;
	wire branch_7_in1_valid;
	wire [0 : 0]branch_7_in2_data;
	wire branch_7_in2_ready;
	wire branch_7_in2_valid;
	wire [0 : 0]branch_7_out1_data;
	wire branch_7_out1_ready;
	wire branch_7_out1_valid;
	wire [0 : 0]branch_7_out2_data;
	wire branch_7_out2_ready;
	wire branch_7_out2_valid;

	wire branch_8_clk;
	wire branch_8_rst;
	wire [31 : 0]branch_8_in1_data;
	wire branch_8_in1_ready;
	wire branch_8_in1_valid;
	wire [0 : 0]branch_8_in2_data;
	wire branch_8_in2_ready;
	wire branch_8_in2_valid;
	wire [31 : 0]branch_8_out1_data;
	wire branch_8_out1_ready;
	wire branch_8_out1_valid;
	wire [31 : 0]branch_8_out2_data;
	wire branch_8_out2_ready;
	wire branch_8_out2_valid;

	wire branch_9_clk;
	wire branch_9_rst;
	wire [2 : 0]branch_9_in1_data;
	wire branch_9_in1_ready;
	wire branch_9_in1_valid;
	wire [0 : 0]branch_9_in2_data;
	wire branch_9_in2_ready;
	wire branch_9_in2_valid;
	wire [2 : 0]branch_9_out1_data;
	wire branch_9_out1_ready;
	wire branch_9_out1_valid;
	wire [2 : 0]branch_9_out2_data;
	wire branch_9_out2_ready;
	wire branch_9_out2_valid;

	wire branch_10_clk;
	wire branch_10_rst;
	wire [4 : 0]branch_10_in1_data;
	wire branch_10_in1_ready;
	wire branch_10_in1_valid;
	wire [0 : 0]branch_10_in2_data;
	wire branch_10_in2_ready;
	wire branch_10_in2_valid;
	wire [4 : 0]branch_10_out1_data;
	wire branch_10_out1_ready;
	wire branch_10_out1_valid;
	wire [4 : 0]branch_10_out2_data;
	wire branch_10_out2_ready;
	wire branch_10_out2_valid;

	wire branch_11_clk;
	wire branch_11_rst;
	wire [4 : 0]branch_11_in1_data;
	wire branch_11_in1_ready;
	wire branch_11_in1_valid;
	wire [0 : 0]branch_11_in2_data;
	wire branch_11_in2_ready;
	wire branch_11_in2_valid;
	wire [4 : 0]branch_11_out1_data;
	wire branch_11_out1_ready;
	wire branch_11_out1_valid;
	wire [4 : 0]branch_11_out2_data;
	wire branch_11_out2_ready;
	wire branch_11_out2_valid;

	wire fork_18_clk;
	wire fork_18_rst;
	wire [0 : 0]fork_18_in1_data;
	wire fork_18_in1_ready;
	wire fork_18_in1_valid;
	wire [0 : 0]fork_18_out1_data;
	wire fork_18_out1_ready;
	wire fork_18_out1_valid;
	wire [0 : 0]fork_18_out2_data;
	wire fork_18_out2_ready;
	wire fork_18_out2_valid;
	wire [0 : 0]fork_18_out3_data;
	wire fork_18_out3_ready;
	wire fork_18_out3_valid;
	wire [0 : 0]fork_18_out4_data;
	wire fork_18_out4_ready;
	wire fork_18_out4_valid;
	wire [0 : 0]fork_18_out5_data;
	wire fork_18_out5_ready;
	wire fork_18_out5_valid;
	wire [0 : 0]fork_18_out6_data;
	wire fork_18_out6_ready;
	wire fork_18_out6_valid;

	wire phiC_18_clk;
	wire phiC_18_rst;
	wire [0 : 0]phiC_18_in1_data;
	wire phiC_18_in1_ready;
	wire phiC_18_in1_valid;
	wire [0 : 0]phiC_18_in2_data;
	wire phiC_18_in2_ready;
	wire phiC_18_in2_valid;
	wire [0 : 0]phiC_18_out1_data;
	wire phiC_18_out1_ready;
	wire phiC_18_out1_valid;
	wire [0 : 0]phiC_18_out2_data;
	wire phiC_18_out2_ready;
	wire phiC_18_out2_valid;

	wire forkC_28_clk;
	wire forkC_28_rst;
	wire [0 : 0]forkC_28_in1_data;
	wire forkC_28_in1_ready;
	wire forkC_28_in1_valid;
	wire [0 : 0]forkC_28_out1_data;
	wire forkC_28_out1_ready;
	wire forkC_28_out1_valid;
	wire [0 : 0]forkC_28_out2_data;
	wire forkC_28_out2_ready;
	wire forkC_28_out2_valid;
	wire [0 : 0]forkC_28_out3_data;
	wire forkC_28_out3_ready;
	wire forkC_28_out3_valid;

	wire branchC_29_clk;
	wire branchC_29_rst;
	wire [0 : 0]branchC_29_in1_data;
	wire branchC_29_in1_ready;
	wire branchC_29_in1_valid;
	wire [0 : 0]branchC_29_in2_data;
	wire branchC_29_in2_ready;
	wire branchC_29_in2_valid;
	wire [0 : 0]branchC_29_out1_data;
	wire branchC_29_out1_ready;
	wire branchC_29_out1_valid;
	wire [0 : 0]branchC_29_out2_data;
	wire branchC_29_out2_ready;
	wire branchC_29_out2_valid;

	wire fork_36_clk;
	wire fork_36_rst;
	wire [0 : 0]fork_36_in1_data;
	wire fork_36_in1_ready;
	wire fork_36_in1_valid;
	wire [0 : 0]fork_36_out1_data;
	wire fork_36_out1_ready;
	wire fork_36_out1_valid;
	wire [0 : 0]fork_36_out2_data;
	wire fork_36_out2_ready;
	wire fork_36_out2_valid;

	wire cst_9_clk;
	wire cst_9_rst;
	wire [0 : 0]cst_9_in1_data;
	wire cst_9_in1_ready;
	wire cst_9_in1_valid;
	wire [0 : 0]cst_9_out1_data;
	wire cst_9_out1_ready;
	wire cst_9_out1_valid;

	wire add_27_clk;
	wire add_27_rst;
	wire [2 : 0]add_27_in1_data;
	wire add_27_in1_ready;
	wire add_27_in1_valid;
	wire [2 : 0]add_27_in2_data;
	wire add_27_in2_ready;
	wire add_27_in2_valid;
	wire [2 : 0]add_27_out1_data;
	wire add_27_out1_ready;
	wire add_27_out1_valid;

	wire cst_10_clk;
	wire cst_10_rst;
	wire [1 : 0]cst_10_in1_data;
	wire cst_10_in1_ready;
	wire cst_10_in1_valid;
	wire [1 : 0]cst_10_out1_data;
	wire cst_10_out1_ready;
	wire cst_10_out1_valid;

	wire icmp_28_clk;
	wire icmp_28_rst;
	wire [2 : 0]icmp_28_in1_data;
	wire icmp_28_in1_ready;
	wire icmp_28_in1_valid;
	wire [2 : 0]icmp_28_in2_data;
	wire icmp_28_in2_ready;
	wire icmp_28_in2_valid;
	wire [0 : 0]icmp_28_out1_data;
	wire icmp_28_out1_ready;
	wire icmp_28_out1_valid;

	wire phi_n8_clk;
	wire phi_n8_rst;
	wire [2 : 0]phi_n8_in1_data;
	wire phi_n8_in1_ready;
	wire phi_n8_in1_valid;
	wire [2 : 0]phi_n8_out1_data;
	wire phi_n8_out1_ready;
	wire phi_n8_out1_valid;

	wire phi_n9_clk;
	wire phi_n9_rst;
	wire [31 : 0]phi_n9_in1_data;
	wire phi_n9_in1_ready;
	wire phi_n9_in1_valid;
	wire [31 : 0]phi_n9_out1_data;
	wire phi_n9_out1_ready;
	wire phi_n9_out1_valid;

	wire phi_n10_clk;
	wire phi_n10_rst;
	wire [4 : 0]phi_n10_in1_data;
	wire phi_n10_in1_ready;
	wire phi_n10_in1_valid;
	wire [4 : 0]phi_n10_out1_data;
	wire phi_n10_out1_ready;
	wire phi_n10_out1_valid;

	wire phi_n11_clk;
	wire phi_n11_rst;
	wire [4 : 0]phi_n11_in1_data;
	wire phi_n11_in1_ready;
	wire phi_n11_in1_valid;
	wire [4 : 0]phi_n11_out1_data;
	wire phi_n11_out1_ready;
	wire phi_n11_out1_valid;

	wire fork_3_clk;
	wire fork_3_rst;
	wire [2 : 0]fork_3_in1_data;
	wire fork_3_in1_ready;
	wire fork_3_in1_valid;
	wire [2 : 0]fork_3_out1_data;
	wire fork_3_out1_ready;
	wire fork_3_out1_valid;
	wire [2 : 0]fork_3_out2_data;
	wire fork_3_out2_ready;
	wire fork_3_out2_valid;

	wire branch_17_clk;
	wire branch_17_rst;
	wire [2 : 0]branch_17_in1_data;
	wire branch_17_in1_ready;
	wire branch_17_in1_valid;
	wire [0 : 0]branch_17_in2_data;
	wire branch_17_in2_ready;
	wire branch_17_in2_valid;
	wire [2 : 0]branch_17_out1_data;
	wire branch_17_out1_ready;
	wire branch_17_out1_valid;
	wire [2 : 0]branch_17_out2_data;
	wire branch_17_out2_ready;
	wire branch_17_out2_valid;

	wire branch_18_clk;
	wire branch_18_rst;
	wire [31 : 0]branch_18_in1_data;
	wire branch_18_in1_ready;
	wire branch_18_in1_valid;
	wire [0 : 0]branch_18_in2_data;
	wire branch_18_in2_ready;
	wire branch_18_in2_valid;
	wire [31 : 0]branch_18_out1_data;
	wire branch_18_out1_ready;
	wire branch_18_out1_valid;
	wire [31 : 0]branch_18_out2_data;
	wire branch_18_out2_ready;
	wire branch_18_out2_valid;

	wire branch_19_clk;
	wire branch_19_rst;
	wire [4 : 0]branch_19_in1_data;
	wire branch_19_in1_ready;
	wire branch_19_in1_valid;
	wire [0 : 0]branch_19_in2_data;
	wire branch_19_in2_ready;
	wire branch_19_in2_valid;
	wire [4 : 0]branch_19_out1_data;
	wire branch_19_out1_ready;
	wire branch_19_out1_valid;
	wire [4 : 0]branch_19_out2_data;
	wire branch_19_out2_ready;
	wire branch_19_out2_valid;

	wire branch_20_clk;
	wire branch_20_rst;
	wire [4 : 0]branch_20_in1_data;
	wire branch_20_in1_ready;
	wire branch_20_in1_valid;
	wire [0 : 0]branch_20_in2_data;
	wire branch_20_in2_ready;
	wire branch_20_in2_valid;
	wire [4 : 0]branch_20_out1_data;
	wire branch_20_out1_ready;
	wire branch_20_out1_valid;
	wire [4 : 0]branch_20_out2_data;
	wire branch_20_out2_ready;
	wire branch_20_out2_valid;

	wire fork_20_clk;
	wire fork_20_rst;
	wire [0 : 0]fork_20_in1_data;
	wire fork_20_in1_ready;
	wire fork_20_in1_valid;
	wire [0 : 0]fork_20_out1_data;
	wire fork_20_out1_ready;
	wire fork_20_out1_valid;
	wire [0 : 0]fork_20_out2_data;
	wire fork_20_out2_ready;
	wire fork_20_out2_valid;
	wire [0 : 0]fork_20_out3_data;
	wire fork_20_out3_ready;
	wire fork_20_out3_valid;
	wire [0 : 0]fork_20_out4_data;
	wire fork_20_out4_ready;
	wire fork_20_out4_valid;
	wire [0 : 0]fork_20_out5_data;
	wire fork_20_out5_ready;
	wire fork_20_out5_valid;

	wire phiC_20_clk;
	wire phiC_20_rst;
	wire [0 : 0]phiC_20_in1_data;
	wire phiC_20_in1_ready;
	wire phiC_20_in1_valid;
	wire [0 : 0]phiC_20_out1_data;
	wire phiC_20_out1_ready;
	wire phiC_20_out1_valid;

	wire branchC_31_clk;
	wire branchC_31_rst;
	wire [0 : 0]branchC_31_in1_data;
	wire branchC_31_in1_ready;
	wire branchC_31_in1_valid;
	wire [0 : 0]branchC_31_in2_data;
	wire branchC_31_in2_ready;
	wire branchC_31_in2_valid;
	wire [0 : 0]branchC_31_out1_data;
	wire branchC_31_out1_ready;
	wire branchC_31_out1_valid;
	wire [0 : 0]branchC_31_out2_data;
	wire branchC_31_out2_ready;
	wire branchC_31_out2_valid;

	wire source_4_clk;
	wire source_4_rst;
	wire [0 : 0]source_4_out1_data;
	wire source_4_out1_ready;
	wire source_4_out1_valid;

	wire source_5_clk;
	wire source_5_rst;
	wire [1 : 0]source_5_out1_data;
	wire source_5_out1_ready;
	wire source_5_out1_valid;

	wire cst_14_clk;
	wire cst_14_rst;
	wire [0 : 0]cst_14_in1_data;
	wire cst_14_in1_ready;
	wire cst_14_in1_valid;
	wire [0 : 0]cst_14_out1_data;
	wire cst_14_out1_ready;
	wire cst_14_out1_valid;

	wire add_37_clk;
	wire add_37_rst;
	wire [4 : 0]add_37_in1_data;
	wire add_37_in1_ready;
	wire add_37_in1_valid;
	wire [4 : 0]add_37_in2_data;
	wire add_37_in2_ready;
	wire add_37_in2_valid;
	wire [4 : 0]add_37_out1_data;
	wire add_37_out1_ready;
	wire add_37_out1_valid;

	wire cst_15_clk;
	wire cst_15_rst;
	wire [4 : 0]cst_15_in1_data;
	wire cst_15_in1_ready;
	wire cst_15_in1_valid;
	wire [4 : 0]cst_15_out1_data;
	wire cst_15_out1_ready;
	wire cst_15_out1_valid;

	wire icmp_38_clk;
	wire icmp_38_rst;
	wire [4 : 0]icmp_38_in1_data;
	wire icmp_38_in1_ready;
	wire icmp_38_in1_valid;
	wire [4 : 0]icmp_38_in2_data;
	wire icmp_38_in2_ready;
	wire icmp_38_in2_valid;
	wire [0 : 0]icmp_38_out1_data;
	wire icmp_38_out1_ready;
	wire icmp_38_out1_valid;

	wire phi_n0_clk;
	wire phi_n0_rst;
	wire [4 : 0]phi_n0_in1_data;
	wire phi_n0_in1_ready;
	wire phi_n0_in1_valid;
	wire [4 : 0]phi_n0_out1_data;
	wire phi_n0_out1_ready;
	wire phi_n0_out1_valid;

	wire phi_n1_clk;
	wire phi_n1_rst;
	wire [31 : 0]phi_n1_in1_data;
	wire phi_n1_in1_ready;
	wire phi_n1_in1_valid;
	wire [31 : 0]phi_n1_out1_data;
	wire phi_n1_out1_ready;
	wire phi_n1_out1_valid;

	wire fork_5_clk;
	wire fork_5_rst;
	wire [4 : 0]fork_5_in1_data;
	wire fork_5_in1_ready;
	wire fork_5_in1_valid;
	wire [4 : 0]fork_5_out1_data;
	wire fork_5_out1_ready;
	wire fork_5_out1_valid;
	wire [4 : 0]fork_5_out2_data;
	wire fork_5_out2_ready;
	wire fork_5_out2_valid;

	wire branch_24_clk;
	wire branch_24_rst;
	wire [31 : 0]branch_24_in1_data;
	wire branch_24_in1_ready;
	wire branch_24_in1_valid;
	wire [0 : 0]branch_24_in2_data;
	wire branch_24_in2_ready;
	wire branch_24_in2_valid;
	wire [31 : 0]branch_24_out1_data;
	wire branch_24_out1_ready;
	wire branch_24_out1_valid;
	wire [31 : 0]branch_24_out2_data;
	wire branch_24_out2_ready;
	wire branch_24_out2_valid;

	wire branch_25_clk;
	wire branch_25_rst;
	wire [4 : 0]branch_25_in1_data;
	wire branch_25_in1_ready;
	wire branch_25_in1_valid;
	wire [0 : 0]branch_25_in2_data;
	wire branch_25_in2_ready;
	wire branch_25_in2_valid;
	wire [4 : 0]branch_25_out1_data;
	wire branch_25_out1_ready;
	wire branch_25_out1_valid;
	wire [4 : 0]branch_25_out2_data;
	wire branch_25_out2_ready;
	wire branch_25_out2_valid;

	wire fork_22_clk;
	wire fork_22_rst;
	wire [0 : 0]fork_22_in1_data;
	wire fork_22_in1_ready;
	wire fork_22_in1_valid;
	wire [0 : 0]fork_22_out1_data;
	wire fork_22_out1_ready;
	wire fork_22_out1_valid;
	wire [0 : 0]fork_22_out2_data;
	wire fork_22_out2_ready;
	wire fork_22_out2_valid;
	wire [0 : 0]fork_22_out3_data;
	wire fork_22_out3_ready;
	wire fork_22_out3_valid;

	wire phiC_22_clk;
	wire phiC_22_rst;
	wire [0 : 0]phiC_22_in1_data;
	wire phiC_22_in1_ready;
	wire phiC_22_in1_valid;
	wire [0 : 0]phiC_22_out1_data;
	wire phiC_22_out1_ready;
	wire phiC_22_out1_valid;

	wire branchC_33_clk;
	wire branchC_33_rst;
	wire [0 : 0]branchC_33_in1_data;
	wire branchC_33_in1_ready;
	wire branchC_33_in1_valid;
	wire [0 : 0]branchC_33_in2_data;
	wire branchC_33_in2_ready;
	wire branchC_33_in2_valid;
	wire [0 : 0]branchC_33_out1_data;
	wire branchC_33_out1_ready;
	wire branchC_33_out1_valid;
	wire [0 : 0]branchC_33_out2_data;
	wire branchC_33_out2_ready;
	wire branchC_33_out2_valid;

	wire source_9_clk;
	wire source_9_rst;
	wire [0 : 0]source_9_out1_data;
	wire source_9_out1_ready;
	wire source_9_out1_valid;

	wire source_10_clk;
	wire source_10_rst;
	wire [4 : 0]source_10_out1_data;
	wire source_10_out1_ready;
	wire source_10_out1_valid;

	wire ret_0_clk;
	wire ret_0_rst;
	wire [31 : 0]ret_0_in1_data;
	wire ret_0_in1_ready;
	wire ret_0_in1_valid;
	wire [31 : 0]ret_0_out1_data;
	wire ret_0_out1_ready;
	wire ret_0_out1_valid;

	wire phi_n15_clk;
	wire phi_n15_rst;
	wire [31 : 0]phi_n15_in1_data;
	wire phi_n15_in1_ready;
	wire phi_n15_in1_valid;
	wire [31 : 0]phi_n15_out1_data;
	wire phi_n15_out1_ready;
	wire phi_n15_out1_valid;

	wire end_0_clk;
	wire end_0_rst;
	wire [0 : 0]end_0_in1_data;
	wire end_0_in1_ready;
	wire end_0_in1_valid;
	wire [0 : 0]end_0_in2_data;
	wire end_0_in2_ready;
	wire end_0_in2_valid;
	wire [0 : 0]end_0_in3_data;
	wire end_0_in3_ready;
	wire end_0_in3_valid;
	wire [31 : 0]end_0_in4_data;
	wire end_0_in4_ready;
	wire end_0_in4_valid;
	wire [31 : 0]end_0_out1_data;
	wire end_0_out1_ready;
	wire end_0_out1_valid;

	wire phiC_23_clk;
	wire phiC_23_rst;
	wire [0 : 0]phiC_23_in1_data;
	wire phiC_23_in1_ready;
	wire phiC_23_in1_valid;
	wire [0 : 0]phiC_23_out1_data;
	wire phiC_23_out1_ready;
	wire phiC_23_out1_valid;

	wire sink_0_clk;
	wire sink_0_rst;
	wire [0 : 0]sink_0_in1_data;
	wire sink_0_in1_ready;
	wire sink_0_in1_valid;

	wire phi_3_clk;
	wire phi_3_rst;
	wire [0 : 0]phi_3_in1_data;
	wire phi_3_in1_ready;
	wire phi_3_in1_valid;
	wire [4 : 0]phi_3_in2_data;
	wire phi_3_in2_ready;
	wire phi_3_in2_valid;
	wire [4 : 0]phi_3_in3_data;
	wire phi_3_in3_ready;
	wire phi_3_in3_valid;
	wire [4 : 0]phi_3_out1_data;
	wire phi_3_out1_ready;
	wire phi_3_out1_valid;

	wire brCst_block3_clk;
	wire brCst_block3_rst;
	wire [0 : 0]brCst_block3_in1_data;
	wire brCst_block3_in1_ready;
	wire brCst_block3_in1_valid;
	wire [0 : 0]brCst_block3_out1_data;
	wire brCst_block3_out1_ready;
	wire brCst_block3_out1_valid;

	wire cst_2_clk;
	wire cst_2_rst;
	wire [0 : 0]cst_2_in1_data;
	wire cst_2_in1_ready;
	wire cst_2_in1_valid;
	wire [0 : 0]cst_2_out1_data;
	wire cst_2_out1_ready;
	wire cst_2_out1_valid;

	wire cst_3_clk;
	wire cst_3_rst;
	wire [0 : 0]cst_3_in1_data;
	wire cst_3_in1_ready;
	wire cst_3_in1_valid;
	wire [0 : 0]cst_3_out1_data;
	wire cst_3_out1_ready;
	wire cst_3_out1_valid;

	wire phi_n2_clk;
	wire phi_n2_rst;
	wire [4 : 0]phi_n2_in1_data;
	wire phi_n2_in1_ready;
	wire phi_n2_in1_valid;
	wire [4 : 0]phi_n2_in2_data;
	wire phi_n2_in2_ready;
	wire phi_n2_in2_valid;
	wire [4 : 0]phi_n2_out1_data;
	wire phi_n2_out1_ready;
	wire phi_n2_out1_valid;

	wire branch_3_clk;
	wire branch_3_rst;
	wire [0 : 0]branch_3_in1_data;
	wire branch_3_in1_ready;
	wire branch_3_in1_valid;
	wire [0 : 0]branch_3_in2_data;
	wire branch_3_in2_ready;
	wire branch_3_in2_valid;
	wire [0 : 0]branch_3_out1_data;
	wire branch_3_out1_ready;
	wire branch_3_out1_valid;
	wire [0 : 0]branch_3_out2_data;
	wire branch_3_out2_ready;
	wire branch_3_out2_valid;

	wire branch_4_clk;
	wire branch_4_rst;
	wire [0 : 0]branch_4_in1_data;
	wire branch_4_in1_ready;
	wire branch_4_in1_valid;
	wire [0 : 0]branch_4_in2_data;
	wire branch_4_in2_ready;
	wire branch_4_in2_valid;
	wire [0 : 0]branch_4_out1_data;
	wire branch_4_out1_ready;
	wire branch_4_out1_valid;
	wire [0 : 0]branch_4_out2_data;
	wire branch_4_out2_ready;
	wire branch_4_out2_valid;

	wire branch_5_clk;
	wire branch_5_rst;
	wire [4 : 0]branch_5_in1_data;
	wire branch_5_in1_ready;
	wire branch_5_in1_valid;
	wire [0 : 0]branch_5_in2_data;
	wire branch_5_in2_ready;
	wire branch_5_in2_valid;
	wire [4 : 0]branch_5_out1_data;
	wire branch_5_out1_ready;
	wire branch_5_out1_valid;
	wire [4 : 0]branch_5_out2_data;
	wire branch_5_out2_ready;
	wire branch_5_out2_valid;

	wire branch_6_clk;
	wire branch_6_rst;
	wire [4 : 0]branch_6_in1_data;
	wire branch_6_in1_ready;
	wire branch_6_in1_valid;
	wire [0 : 0]branch_6_in2_data;
	wire branch_6_in2_ready;
	wire branch_6_in2_valid;
	wire [4 : 0]branch_6_out1_data;
	wire branch_6_out1_ready;
	wire branch_6_out1_valid;
	wire [4 : 0]branch_6_out2_data;
	wire branch_6_out2_ready;
	wire branch_6_out2_valid;

	wire fork_17_clk;
	wire fork_17_rst;
	wire [0 : 0]fork_17_in1_data;
	wire fork_17_in1_ready;
	wire fork_17_in1_valid;
	wire [0 : 0]fork_17_out1_data;
	wire fork_17_out1_ready;
	wire fork_17_out1_valid;
	wire [0 : 0]fork_17_out2_data;
	wire fork_17_out2_ready;
	wire fork_17_out2_valid;
	wire [0 : 0]fork_17_out3_data;
	wire fork_17_out3_ready;
	wire fork_17_out3_valid;
	wire [0 : 0]fork_17_out4_data;
	wire fork_17_out4_ready;
	wire fork_17_out4_valid;
	wire [0 : 0]fork_17_out5_data;
	wire fork_17_out5_ready;
	wire fork_17_out5_valid;

	wire phiC_17_clk;
	wire phiC_17_rst;
	wire [0 : 0]phiC_17_in1_data;
	wire phiC_17_in1_ready;
	wire phiC_17_in1_valid;
	wire [0 : 0]phiC_17_in2_data;
	wire phiC_17_in2_ready;
	wire phiC_17_in2_valid;
	wire [0 : 0]phiC_17_out1_data;
	wire phiC_17_out1_ready;
	wire phiC_17_out1_valid;
	wire [0 : 0]phiC_17_out2_data;
	wire phiC_17_out2_ready;
	wire phiC_17_out2_valid;

	wire forkC_27_clk;
	wire forkC_27_rst;
	wire [0 : 0]forkC_27_in1_data;
	wire forkC_27_in1_ready;
	wire forkC_27_in1_valid;
	wire [0 : 0]forkC_27_out1_data;
	wire forkC_27_out1_ready;
	wire forkC_27_out1_valid;
	wire [0 : 0]forkC_27_out2_data;
	wire forkC_27_out2_ready;
	wire forkC_27_out2_valid;
	wire [0 : 0]forkC_27_out3_data;
	wire forkC_27_out3_ready;
	wire forkC_27_out3_valid;
	wire [0 : 0]forkC_27_out4_data;
	wire forkC_27_out4_ready;
	wire forkC_27_out4_valid;

	wire branchC_28_clk;
	wire branchC_28_rst;
	wire [0 : 0]branchC_28_in1_data;
	wire branchC_28_in1_ready;
	wire branchC_28_in1_valid;
	wire [0 : 0]branchC_28_in2_data;
	wire branchC_28_in2_ready;
	wire branchC_28_in2_valid;
	wire [0 : 0]branchC_28_out1_data;
	wire branchC_28_out1_ready;
	wire branchC_28_out1_valid;
	wire [0 : 0]branchC_28_out2_data;
	wire branchC_28_out2_ready;
	wire branchC_28_out2_valid;

	wire cst_11_clk;
	wire cst_11_rst;
	wire [4 : 0]cst_11_in1_data;
	wire cst_11_in1_ready;
	wire cst_11_in1_valid;
	wire [4 : 0]cst_11_out1_data;
	wire cst_11_out1_ready;
	wire cst_11_out1_valid;

	wire mul_30_clk;
	wire mul_30_rst;
	wire [4 : 0]mul_30_in1_data;
	wire mul_30_in1_ready;
	wire mul_30_in1_valid;
	wire [4 : 0]mul_30_in2_data;
	wire mul_30_in2_ready;
	wire mul_30_in2_valid;
	wire [9 : 0]mul_30_out1_data;
	wire mul_30_out1_ready;
	wire mul_30_out1_valid;

	wire add_31_clk;
	wire add_31_rst;
	wire [10 : 0]add_31_in1_data;
	wire add_31_in1_ready;
	wire add_31_in1_valid;
	wire [10 : 0]add_31_in2_data;
	wire add_31_in2_ready;
	wire add_31_in2_valid;
	wire [10 : 0]add_31_out1_data;
	wire add_31_out1_ready;
	wire add_31_out1_valid;

	wire store_0_clk;
	wire store_0_rst;
	wire [31 : 0]store_0_in1_data;
	wire store_0_in1_ready;
	wire store_0_in1_valid;
	wire [10 : 0]store_0_in2_data;
	wire store_0_in2_ready;
	wire store_0_in2_valid;
	wire [31 : 0]store_0_out1_data;
	wire store_0_out1_ready;
	wire store_0_out1_valid;
	wire [10 : 0]store_0_out2_data;
	wire store_0_out2_ready;
	wire store_0_out2_valid;

	wire cst_12_clk;
	wire cst_12_rst;
	wire [0 : 0]cst_12_in1_data;
	wire cst_12_in1_ready;
	wire cst_12_in1_valid;
	wire [0 : 0]cst_12_out1_data;
	wire cst_12_out1_ready;
	wire cst_12_out1_valid;

	wire add_34_clk;
	wire add_34_rst;
	wire [4 : 0]add_34_in1_data;
	wire add_34_in1_ready;
	wire add_34_in1_valid;
	wire [4 : 0]add_34_in2_data;
	wire add_34_in2_ready;
	wire add_34_in2_valid;
	wire [4 : 0]add_34_out1_data;
	wire add_34_out1_ready;
	wire add_34_out1_valid;

	wire cst_13_clk;
	wire cst_13_rst;
	wire [4 : 0]cst_13_in1_data;
	wire cst_13_in1_ready;
	wire cst_13_in1_valid;
	wire [4 : 0]cst_13_out1_data;
	wire cst_13_out1_ready;
	wire cst_13_out1_valid;

	wire icmp_35_clk;
	wire icmp_35_rst;
	wire [4 : 0]icmp_35_in1_data;
	wire icmp_35_in1_ready;
	wire icmp_35_in1_valid;
	wire [4 : 0]icmp_35_in2_data;
	wire icmp_35_in2_ready;
	wire icmp_35_in2_valid;
	wire [0 : 0]icmp_35_out1_data;
	wire icmp_35_out1_ready;
	wire icmp_35_out1_valid;

	wire phi_n3_clk;
	wire phi_n3_rst;
	wire [4 : 0]phi_n3_in1_data;
	wire phi_n3_in1_ready;
	wire phi_n3_in1_valid;
	wire [4 : 0]phi_n3_out1_data;
	wire phi_n3_out1_ready;
	wire phi_n3_out1_valid;

	wire phi_n4_clk;
	wire phi_n4_rst;
	wire [4 : 0]phi_n4_in1_data;
	wire phi_n4_in1_ready;
	wire phi_n4_in1_valid;
	wire [4 : 0]phi_n4_out1_data;
	wire phi_n4_out1_ready;
	wire phi_n4_out1_valid;

	wire phi_n5_clk;
	wire phi_n5_rst;
	wire [31 : 0]phi_n5_in1_data;
	wire phi_n5_in1_ready;
	wire phi_n5_in1_valid;
	wire [31 : 0]phi_n5_out1_data;
	wire phi_n5_out1_ready;
	wire phi_n5_out1_valid;

	wire fork_4_clk;
	wire fork_4_rst;
	wire [4 : 0]fork_4_in1_data;
	wire fork_4_in1_ready;
	wire fork_4_in1_valid;
	wire [4 : 0]fork_4_out1_data;
	wire fork_4_out1_ready;
	wire fork_4_out1_valid;
	wire [4 : 0]fork_4_out2_data;
	wire fork_4_out2_ready;
	wire fork_4_out2_valid;

	wire fork_6_clk;
	wire fork_6_rst;
	wire [4 : 0]fork_6_in1_data;
	wire fork_6_in1_ready;
	wire fork_6_in1_valid;
	wire [4 : 0]fork_6_out1_data;
	wire fork_6_out1_ready;
	wire fork_6_out1_valid;
	wire [4 : 0]fork_6_out2_data;
	wire fork_6_out2_ready;
	wire fork_6_out2_valid;

	wire fork_7_clk;
	wire fork_7_rst;
	wire [4 : 0]fork_7_in1_data;
	wire fork_7_in1_ready;
	wire fork_7_in1_valid;
	wire [4 : 0]fork_7_out1_data;
	wire fork_7_out1_ready;
	wire fork_7_out1_valid;
	wire [4 : 0]fork_7_out2_data;
	wire fork_7_out2_ready;
	wire fork_7_out2_valid;

	wire fork_8_clk;
	wire fork_8_rst;
	wire [31 : 0]fork_8_in1_data;
	wire fork_8_in1_ready;
	wire fork_8_in1_valid;
	wire [31 : 0]fork_8_out1_data;
	wire fork_8_out1_ready;
	wire fork_8_out1_valid;
	wire [31 : 0]fork_8_out2_data;
	wire fork_8_out2_ready;
	wire fork_8_out2_valid;

	wire branch_21_clk;
	wire branch_21_rst;
	wire [4 : 0]branch_21_in1_data;
	wire branch_21_in1_ready;
	wire branch_21_in1_valid;
	wire [0 : 0]branch_21_in2_data;
	wire branch_21_in2_ready;
	wire branch_21_in2_valid;
	wire [4 : 0]branch_21_out1_data;
	wire branch_21_out1_ready;
	wire branch_21_out1_valid;
	wire [4 : 0]branch_21_out2_data;
	wire branch_21_out2_ready;
	wire branch_21_out2_valid;

	wire branch_22_clk;
	wire branch_22_rst;
	wire [4 : 0]branch_22_in1_data;
	wire branch_22_in1_ready;
	wire branch_22_in1_valid;
	wire [0 : 0]branch_22_in2_data;
	wire branch_22_in2_ready;
	wire branch_22_in2_valid;
	wire [4 : 0]branch_22_out1_data;
	wire branch_22_out1_ready;
	wire branch_22_out1_valid;
	wire [4 : 0]branch_22_out2_data;
	wire branch_22_out2_ready;
	wire branch_22_out2_valid;

	wire branch_23_clk;
	wire branch_23_rst;
	wire [31 : 0]branch_23_in1_data;
	wire branch_23_in1_ready;
	wire branch_23_in1_valid;
	wire [0 : 0]branch_23_in2_data;
	wire branch_23_in2_ready;
	wire branch_23_in2_valid;
	wire [31 : 0]branch_23_out1_data;
	wire branch_23_out1_ready;
	wire branch_23_out1_valid;
	wire [31 : 0]branch_23_out2_data;
	wire branch_23_out2_ready;
	wire branch_23_out2_valid;

	wire fork_21_clk;
	wire fork_21_rst;
	wire [0 : 0]fork_21_in1_data;
	wire fork_21_in1_ready;
	wire fork_21_in1_valid;
	wire [0 : 0]fork_21_out1_data;
	wire fork_21_out1_ready;
	wire fork_21_out1_valid;
	wire [0 : 0]fork_21_out2_data;
	wire fork_21_out2_ready;
	wire fork_21_out2_valid;
	wire [0 : 0]fork_21_out3_data;
	wire fork_21_out3_ready;
	wire fork_21_out3_valid;
	wire [0 : 0]fork_21_out4_data;
	wire fork_21_out4_ready;
	wire fork_21_out4_valid;

	wire cst_16_clk;
	wire cst_16_rst;
	wire [0 : 0]cst_16_in1_data;
	wire cst_16_in1_ready;
	wire cst_16_in1_valid;
	wire [0 : 0]cst_16_out1_data;
	wire cst_16_out1_ready;
	wire cst_16_out1_valid;

	wire phiC_21_clk;
	wire phiC_21_rst;
	wire [0 : 0]phiC_21_in1_data;
	wire phiC_21_in1_ready;
	wire phiC_21_in1_valid;
	wire [0 : 0]phiC_21_out1_data;
	wire phiC_21_out1_ready;
	wire phiC_21_out1_valid;

	wire forkC_31_clk;
	wire forkC_31_rst;
	wire [0 : 0]forkC_31_in1_data;
	wire forkC_31_in1_ready;
	wire forkC_31_in1_valid;
	wire [0 : 0]forkC_31_out1_data;
	wire forkC_31_out1_ready;
	wire forkC_31_out1_valid;
	wire [0 : 0]forkC_31_out2_data;
	wire forkC_31_out2_ready;
	wire forkC_31_out2_valid;

	wire branchC_32_clk;
	wire branchC_32_rst;
	wire [0 : 0]branchC_32_in1_data;
	wire branchC_32_in1_ready;
	wire branchC_32_in1_valid;
	wire [0 : 0]branchC_32_in2_data;
	wire branchC_32_in2_ready;
	wire branchC_32_in2_valid;
	wire [0 : 0]branchC_32_out1_data;
	wire branchC_32_out1_ready;
	wire branchC_32_out1_valid;
	wire [0 : 0]branchC_32_out2_data;
	wire branchC_32_out2_ready;
	wire branchC_32_out2_valid;

	wire source_6_clk;
	wire source_6_rst;
	wire [4 : 0]source_6_out1_data;
	wire source_6_out1_ready;
	wire source_6_out1_valid;

	wire source_7_clk;
	wire source_7_rst;
	wire [0 : 0]source_7_out1_data;
	wire source_7_out1_ready;
	wire source_7_out1_valid;

	wire source_8_clk;
	wire source_8_rst;
	wire [4 : 0]source_8_out1_data;
	wire source_8_out1_ready;
	wire source_8_out1_valid;

	wire phi_1_clk;
	wire phi_1_rst;
	wire [0 : 0]phi_1_in1_data;
	wire phi_1_in1_ready;
	wire phi_1_in1_valid;
	wire [4 : 0]phi_1_in2_data;
	wire phi_1_in2_ready;
	wire phi_1_in2_valid;
	wire [4 : 0]phi_1_in3_data;
	wire phi_1_in3_ready;
	wire phi_1_in3_valid;
	wire [4 : 0]phi_1_out1_data;
	wire phi_1_out1_ready;
	wire phi_1_out1_valid;

	wire brCst_block2_clk;
	wire brCst_block2_rst;
	wire [0 : 0]brCst_block2_in1_data;
	wire brCst_block2_in1_ready;
	wire brCst_block2_in1_valid;
	wire [0 : 0]brCst_block2_out1_data;
	wire brCst_block2_out1_ready;
	wire brCst_block2_out1_valid;

	wire cst_1_clk;
	wire cst_1_rst;
	wire [0 : 0]cst_1_in1_data;
	wire cst_1_in1_ready;
	wire cst_1_in1_valid;
	wire [0 : 0]cst_1_out1_data;
	wire cst_1_out1_ready;
	wire cst_1_out1_valid;

	wire branch_1_clk;
	wire branch_1_rst;
	wire [0 : 0]branch_1_in1_data;
	wire branch_1_in1_ready;
	wire branch_1_in1_valid;
	wire [0 : 0]branch_1_in2_data;
	wire branch_1_in2_ready;
	wire branch_1_in2_valid;
	wire [0 : 0]branch_1_out1_data;
	wire branch_1_out1_ready;
	wire branch_1_out1_valid;
	wire [0 : 0]branch_1_out2_data;
	wire branch_1_out2_ready;
	wire branch_1_out2_valid;

	wire branch_2_clk;
	wire branch_2_rst;
	wire [4 : 0]branch_2_in1_data;
	wire branch_2_in1_ready;
	wire branch_2_in1_valid;
	wire [0 : 0]branch_2_in2_data;
	wire branch_2_in2_ready;
	wire branch_2_in2_valid;
	wire [4 : 0]branch_2_out1_data;
	wire branch_2_out1_ready;
	wire branch_2_out1_valid;
	wire [4 : 0]branch_2_out2_data;
	wire branch_2_out2_ready;
	wire branch_2_out2_valid;

	wire fork_16_clk;
	wire fork_16_rst;
	wire [0 : 0]fork_16_in1_data;
	wire fork_16_in1_ready;
	wire fork_16_in1_valid;
	wire [0 : 0]fork_16_out1_data;
	wire fork_16_out1_ready;
	wire fork_16_out1_valid;
	wire [0 : 0]fork_16_out2_data;
	wire fork_16_out2_ready;
	wire fork_16_out2_valid;
	wire [0 : 0]fork_16_out3_data;
	wire fork_16_out3_ready;
	wire fork_16_out3_valid;

	wire phiC_16_clk;
	wire phiC_16_rst;
	wire [0 : 0]phiC_16_in1_data;
	wire phiC_16_in1_ready;
	wire phiC_16_in1_valid;
	wire [0 : 0]phiC_16_in2_data;
	wire phiC_16_in2_ready;
	wire phiC_16_in2_valid;
	wire [0 : 0]phiC_16_out1_data;
	wire phiC_16_out1_ready;
	wire phiC_16_out1_valid;
	wire [0 : 0]phiC_16_out2_data;
	wire phiC_16_out2_ready;
	wire phiC_16_out2_valid;

	wire forkC_26_clk;
	wire forkC_26_rst;
	wire [0 : 0]forkC_26_in1_data;
	wire forkC_26_in1_ready;
	wire forkC_26_in1_valid;
	wire [0 : 0]forkC_26_out1_data;
	wire forkC_26_out1_ready;
	wire forkC_26_out1_valid;
	wire [0 : 0]forkC_26_out2_data;
	wire forkC_26_out2_ready;
	wire forkC_26_out2_valid;
	wire [0 : 0]forkC_26_out3_data;
	wire forkC_26_out3_ready;
	wire forkC_26_out3_valid;

	wire branchC_27_clk;
	wire branchC_27_rst;
	wire [0 : 0]branchC_27_in1_data;
	wire branchC_27_in1_ready;
	wire branchC_27_in1_valid;
	wire [0 : 0]branchC_27_in2_data;
	wire branchC_27_in2_ready;
	wire branchC_27_in2_valid;
	wire [0 : 0]branchC_27_out1_data;
	wire branchC_27_out1_ready;
	wire branchC_27_out1_valid;
	wire [0 : 0]branchC_27_out2_data;
	wire branchC_27_out2_ready;
	wire branchC_27_out2_valid;

	wire phi_8_clk;
	wire phi_8_rst;
	wire [0 : 0]phi_8_in1_data;
	wire phi_8_in1_ready;
	wire phi_8_in1_valid;
	wire [2 : 0]phi_8_in2_data;
	wire phi_8_in2_ready;
	wire phi_8_in2_valid;
	wire [2 : 0]phi_8_in3_data;
	wire phi_8_in3_ready;
	wire phi_8_in3_valid;
	wire [2 : 0]phi_8_out1_data;
	wire phi_8_out1_ready;
	wire phi_8_out1_valid;

	wire phi_9_clk;
	wire phi_9_rst;
	wire [0 : 0]phi_9_in1_data;
	wire phi_9_in1_ready;
	wire phi_9_in1_valid;
	wire [31 : 0]phi_9_in2_data;
	wire phi_9_in2_ready;
	wire phi_9_in2_valid;
	wire [31 : 0]phi_9_in3_data;
	wire phi_9_in3_ready;
	wire phi_9_in3_valid;
	wire [31 : 0]phi_9_out1_data;
	wire phi_9_out1_ready;
	wire phi_9_out1_valid;

	wire cst_5_clk;
	wire cst_5_rst;
	wire [1 : 0]cst_5_in1_data;
	wire cst_5_in1_ready;
	wire cst_5_in1_valid;
	wire [1 : 0]cst_5_out1_data;
	wire cst_5_out1_ready;
	wire cst_5_out1_valid;

	wire mul_10_clk;
	wire mul_10_rst;
	wire [1 : 0]mul_10_in1_data;
	wire mul_10_in1_ready;
	wire mul_10_in1_valid;
	wire [2 : 0]mul_10_in2_data;
	wire mul_10_in2_ready;
	wire mul_10_in2_valid;
	wire [4 : 0]mul_10_out1_data;
	wire mul_10_out1_ready;
	wire mul_10_out1_valid;

	wire add_11_clk;
	wire add_11_rst;
	wire [5 : 0]add_11_in1_data;
	wire add_11_in1_ready;
	wire add_11_in1_valid;
	wire [5 : 0]add_11_in2_data;
	wire add_11_in2_ready;
	wire add_11_in2_valid;
	wire [5 : 0]add_11_out1_data;
	wire add_11_out1_ready;
	wire add_11_out1_valid;

	wire load_14_clk;
	wire load_14_rst;
	wire [31 : 0]load_14_in1_data;
	wire load_14_in1_ready;
	wire load_14_in1_valid;
	wire [5 : 0]load_14_in2_data;
	wire load_14_in2_ready;
	wire load_14_in2_valid;
	wire [31 : 0]load_14_out1_data;
	wire load_14_out1_ready;
	wire load_14_out1_valid;
	wire [5 : 0]load_14_out2_data;
	wire load_14_out2_ready;
	wire load_14_out2_valid;

	wire add_15_clk;
	wire add_15_rst;
	wire [5 : 0]add_15_in1_data;
	wire add_15_in1_ready;
	wire add_15_in1_valid;
	wire [5 : 0]add_15_in2_data;
	wire add_15_in2_ready;
	wire add_15_in2_valid;
	wire [5 : 0]add_15_out1_data;
	wire add_15_out1_ready;
	wire add_15_out1_valid;

	wire cst_6_clk;
	wire cst_6_rst;
	wire [4 : 0]cst_6_in1_data;
	wire cst_6_in1_ready;
	wire cst_6_in1_valid;
	wire [4 : 0]cst_6_out1_data;
	wire cst_6_out1_ready;
	wire cst_6_out1_valid;

	wire mul_16_clk;
	wire mul_16_rst;
	wire [4 : 0]mul_16_in1_data;
	wire mul_16_in1_ready;
	wire mul_16_in1_valid;
	wire [5 : 0]mul_16_in2_data;
	wire mul_16_in2_ready;
	wire mul_16_in2_valid;
	wire [10 : 0]mul_16_out1_data;
	wire mul_16_out1_ready;
	wire mul_16_out1_valid;

	wire add_17_clk;
	wire add_17_rst;
	wire [11 : 0]add_17_in1_data;
	wire add_17_in1_ready;
	wire add_17_in1_valid;
	wire [11 : 0]add_17_in2_data;
	wire add_17_in2_ready;
	wire add_17_in2_valid;
	wire [11 : 0]add_17_out1_data;
	wire add_17_out1_ready;
	wire add_17_out1_valid;

	wire add_18_clk;
	wire add_18_rst;
	wire [12 : 0]add_18_in1_data;
	wire add_18_in1_ready;
	wire add_18_in1_valid;
	wire [12 : 0]add_18_in2_data;
	wire add_18_in2_ready;
	wire add_18_in2_valid;
	wire [12 : 0]add_18_out1_data;
	wire add_18_out1_ready;
	wire add_18_out1_valid;

	wire load_21_clk;
	wire load_21_rst;
	wire [31 : 0]load_21_in1_data;
	wire load_21_in1_ready;
	wire load_21_in1_valid;
	wire [12 : 0]load_21_in2_data;
	wire load_21_in2_ready;
	wire load_21_in2_valid;
	wire [31 : 0]load_21_out1_data;
	wire load_21_out1_ready;
	wire load_21_out1_valid;
	wire [12 : 0]load_21_out2_data;
	wire load_21_out2_ready;
	wire load_21_out2_valid;

	wire mul_22_clk;
	wire mul_22_rst;
	wire [15 : 0]mul_22_in1_data;
	wire mul_22_in1_ready;
	wire mul_22_in1_valid;
	wire [15 : 0]mul_22_in2_data;
	wire mul_22_in2_ready;
	wire mul_22_in2_valid;
	wire [31 : 0]mul_22_out1_data;
	wire mul_22_out1_ready;
	wire mul_22_out1_valid;

	wire add_23_clk;
	wire add_23_rst;
	wire [31 : 0]add_23_in1_data;
	wire add_23_in1_ready;
	wire add_23_in1_valid;
	wire [31 : 0]add_23_in2_data;
	wire add_23_in2_ready;
	wire add_23_in2_valid;
	wire [31 : 0]add_23_out1_data;
	wire add_23_out1_ready;
	wire add_23_out1_valid;

	wire cst_7_clk;
	wire cst_7_rst;
	wire [0 : 0]cst_7_in1_data;
	wire cst_7_in1_ready;
	wire cst_7_in1_valid;
	wire [0 : 0]cst_7_out1_data;
	wire cst_7_out1_ready;
	wire cst_7_out1_valid;

	wire add_24_clk;
	wire add_24_rst;
	wire [2 : 0]add_24_in1_data;
	wire add_24_in1_ready;
	wire add_24_in1_valid;
	wire [2 : 0]add_24_in2_data;
	wire add_24_in2_ready;
	wire add_24_in2_valid;
	wire [2 : 0]add_24_out1_data;
	wire add_24_out1_ready;
	wire add_24_out1_valid;

	wire cst_8_clk;
	wire cst_8_rst;
	wire [1 : 0]cst_8_in1_data;
	wire cst_8_in1_ready;
	wire cst_8_in1_valid;
	wire [1 : 0]cst_8_out1_data;
	wire cst_8_out1_ready;
	wire cst_8_out1_valid;

	wire icmp_25_clk;
	wire icmp_25_rst;
	wire [2 : 0]icmp_25_in1_data;
	wire icmp_25_in1_ready;
	wire icmp_25_in1_valid;
	wire [2 : 0]icmp_25_in2_data;
	wire icmp_25_in2_ready;
	wire icmp_25_in2_valid;
	wire [0 : 0]icmp_25_out1_data;
	wire icmp_25_out1_ready;
	wire icmp_25_out1_valid;

	wire phi_n12_clk;
	wire phi_n12_rst;
	wire [2 : 0]phi_n12_in1_data;
	wire phi_n12_in1_ready;
	wire phi_n12_in1_valid;
	wire [2 : 0]phi_n12_in2_data;
	wire phi_n12_in2_ready;
	wire phi_n12_in2_valid;
	wire [2 : 0]phi_n12_out1_data;
	wire phi_n12_out1_ready;
	wire phi_n12_out1_valid;

	wire phi_n13_clk;
	wire phi_n13_rst;
	wire [4 : 0]phi_n13_in1_data;
	wire phi_n13_in1_ready;
	wire phi_n13_in1_valid;
	wire [4 : 0]phi_n13_in2_data;
	wire phi_n13_in2_ready;
	wire phi_n13_in2_valid;
	wire [4 : 0]phi_n13_out1_data;
	wire phi_n13_out1_ready;
	wire phi_n13_out1_valid;

	wire phi_n14_clk;
	wire phi_n14_rst;
	wire [4 : 0]phi_n14_in1_data;
	wire phi_n14_in1_ready;
	wire phi_n14_in1_valid;
	wire [4 : 0]phi_n14_in2_data;
	wire phi_n14_in2_ready;
	wire phi_n14_in2_valid;
	wire [4 : 0]phi_n14_out1_data;
	wire phi_n14_out1_ready;
	wire phi_n14_out1_valid;

	wire fork_0_clk;
	wire fork_0_rst;
	wire [2 : 0]fork_0_in1_data;
	wire fork_0_in1_ready;
	wire fork_0_in1_valid;
	wire [2 : 0]fork_0_out1_data;
	wire fork_0_out1_ready;
	wire fork_0_out1_valid;
	wire [2 : 0]fork_0_out2_data;
	wire fork_0_out2_ready;
	wire fork_0_out2_valid;
	wire [2 : 0]fork_0_out3_data;
	wire fork_0_out3_ready;
	wire fork_0_out3_valid;

	wire fork_2_clk;
	wire fork_2_rst;
	wire [2 : 0]fork_2_in1_data;
	wire fork_2_in1_ready;
	wire fork_2_in1_valid;
	wire [2 : 0]fork_2_out1_data;
	wire fork_2_out1_ready;
	wire fork_2_out1_valid;
	wire [2 : 0]fork_2_out2_data;
	wire fork_2_out2_ready;
	wire fork_2_out2_valid;

	wire fork_12_clk;
	wire fork_12_rst;
	wire [2 : 0]fork_12_in1_data;
	wire fork_12_in1_ready;
	wire fork_12_in1_valid;
	wire [2 : 0]fork_12_out1_data;
	wire fork_12_out1_ready;
	wire fork_12_out1_valid;
	wire [2 : 0]fork_12_out2_data;
	wire fork_12_out2_ready;
	wire fork_12_out2_valid;
	wire [2 : 0]fork_12_out3_data;
	wire fork_12_out3_ready;
	wire fork_12_out3_valid;

	wire fork_13_clk;
	wire fork_13_rst;
	wire [4 : 0]fork_13_in1_data;
	wire fork_13_in1_ready;
	wire fork_13_in1_valid;
	wire [4 : 0]fork_13_out1_data;
	wire fork_13_out1_ready;
	wire fork_13_out1_valid;
	wire [4 : 0]fork_13_out2_data;
	wire fork_13_out2_ready;
	wire fork_13_out2_valid;

	wire fork_14_clk;
	wire fork_14_rst;
	wire [4 : 0]fork_14_in1_data;
	wire fork_14_in1_ready;
	wire fork_14_in1_valid;
	wire [4 : 0]fork_14_out1_data;
	wire fork_14_out1_ready;
	wire fork_14_out1_valid;
	wire [4 : 0]fork_14_out2_data;
	wire fork_14_out2_ready;
	wire fork_14_out2_valid;

	wire branch_12_clk;
	wire branch_12_rst;
	wire [31 : 0]branch_12_in1_data;
	wire branch_12_in1_ready;
	wire branch_12_in1_valid;
	wire [0 : 0]branch_12_in2_data;
	wire branch_12_in2_ready;
	wire branch_12_in2_valid;
	wire [31 : 0]branch_12_out1_data;
	wire branch_12_out1_ready;
	wire branch_12_out1_valid;
	wire [31 : 0]branch_12_out2_data;
	wire branch_12_out2_ready;
	wire branch_12_out2_valid;

	wire branch_13_clk;
	wire branch_13_rst;
	wire [2 : 0]branch_13_in1_data;
	wire branch_13_in1_ready;
	wire branch_13_in1_valid;
	wire [0 : 0]branch_13_in2_data;
	wire branch_13_in2_ready;
	wire branch_13_in2_valid;
	wire [2 : 0]branch_13_out1_data;
	wire branch_13_out1_ready;
	wire branch_13_out1_valid;
	wire [2 : 0]branch_13_out2_data;
	wire branch_13_out2_ready;
	wire branch_13_out2_valid;

	wire branch_14_clk;
	wire branch_14_rst;
	wire [2 : 0]branch_14_in1_data;
	wire branch_14_in1_ready;
	wire branch_14_in1_valid;
	wire [0 : 0]branch_14_in2_data;
	wire branch_14_in2_ready;
	wire branch_14_in2_valid;
	wire [2 : 0]branch_14_out1_data;
	wire branch_14_out1_ready;
	wire branch_14_out1_valid;
	wire [2 : 0]branch_14_out2_data;
	wire branch_14_out2_ready;
	wire branch_14_out2_valid;

	wire branch_15_clk;
	wire branch_15_rst;
	wire [4 : 0]branch_15_in1_data;
	wire branch_15_in1_ready;
	wire branch_15_in1_valid;
	wire [0 : 0]branch_15_in2_data;
	wire branch_15_in2_ready;
	wire branch_15_in2_valid;
	wire [4 : 0]branch_15_out1_data;
	wire branch_15_out1_ready;
	wire branch_15_out1_valid;
	wire [4 : 0]branch_15_out2_data;
	wire branch_15_out2_ready;
	wire branch_15_out2_valid;

	wire branch_16_clk;
	wire branch_16_rst;
	wire [4 : 0]branch_16_in1_data;
	wire branch_16_in1_ready;
	wire branch_16_in1_valid;
	wire [0 : 0]branch_16_in2_data;
	wire branch_16_in2_ready;
	wire branch_16_in2_valid;
	wire [4 : 0]branch_16_out1_data;
	wire branch_16_out1_ready;
	wire branch_16_out1_valid;
	wire [4 : 0]branch_16_out2_data;
	wire branch_16_out2_ready;
	wire branch_16_out2_valid;

	wire fork_19_clk;
	wire fork_19_rst;
	wire [0 : 0]fork_19_in1_data;
	wire fork_19_in1_ready;
	wire fork_19_in1_valid;
	wire [0 : 0]fork_19_out1_data;
	wire fork_19_out1_ready;
	wire fork_19_out1_valid;
	wire [0 : 0]fork_19_out2_data;
	wire fork_19_out2_ready;
	wire fork_19_out2_valid;
	wire [0 : 0]fork_19_out3_data;
	wire fork_19_out3_ready;
	wire fork_19_out3_valid;
	wire [0 : 0]fork_19_out4_data;
	wire fork_19_out4_ready;
	wire fork_19_out4_valid;
	wire [0 : 0]fork_19_out5_data;
	wire fork_19_out5_ready;
	wire fork_19_out5_valid;
	wire [0 : 0]fork_19_out6_data;
	wire fork_19_out6_ready;
	wire fork_19_out6_valid;

	wire phiC_19_clk;
	wire phiC_19_rst;
	wire [0 : 0]phiC_19_in1_data;
	wire phiC_19_in1_ready;
	wire phiC_19_in1_valid;
	wire [0 : 0]phiC_19_in2_data;
	wire phiC_19_in2_ready;
	wire phiC_19_in2_valid;
	wire [0 : 0]phiC_19_out1_data;
	wire phiC_19_out1_ready;
	wire phiC_19_out1_valid;
	wire [0 : 0]phiC_19_out2_data;
	wire phiC_19_out2_ready;
	wire phiC_19_out2_valid;

	wire branchC_30_clk;
	wire branchC_30_rst;
	wire [0 : 0]branchC_30_in1_data;
	wire branchC_30_in1_ready;
	wire branchC_30_in1_valid;
	wire [0 : 0]branchC_30_in2_data;
	wire branchC_30_in2_ready;
	wire branchC_30_in2_valid;
	wire [0 : 0]branchC_30_out1_data;
	wire branchC_30_out1_ready;
	wire branchC_30_out1_valid;
	wire [0 : 0]branchC_30_out2_data;
	wire branchC_30_out2_ready;
	wire branchC_30_out2_valid;

	wire source_0_clk;
	wire source_0_rst;
	wire [1 : 0]source_0_out1_data;
	wire source_0_out1_ready;
	wire source_0_out1_valid;

	wire source_1_clk;
	wire source_1_rst;
	wire [4 : 0]source_1_out1_data;
	wire source_1_out1_ready;
	wire source_1_out1_valid;

	wire source_2_clk;
	wire source_2_rst;
	wire [0 : 0]source_2_out1_data;
	wire source_2_out1_ready;
	wire source_2_out1_valid;

	wire source_3_clk;
	wire source_3_rst;
	wire [1 : 0]source_3_out1_data;
	wire source_3_out1_ready;
	wire source_3_out1_valid;

	wire fork_37_clk;
	wire fork_37_rst;
	wire [0 : 0]fork_37_in1_data;
	wire fork_37_in1_ready;
	wire fork_37_in1_valid;
	wire [0 : 0]fork_37_out1_data;
	wire fork_37_out1_ready;
	wire fork_37_out1_valid;
	wire [0 : 0]fork_37_out2_data;
	wire fork_37_out2_ready;
	wire fork_37_out2_valid;

	wire brCst_block1_clk;
	wire brCst_block1_rst;
	wire [0 : 0]brCst_block1_in1_data;
	wire brCst_block1_in1_ready;
	wire brCst_block1_in1_valid;
	wire [0 : 0]brCst_block1_out1_data;
	wire brCst_block1_out1_ready;
	wire brCst_block1_out1_valid;

	wire cst_0_clk;
	wire cst_0_rst;
	wire [0 : 0]cst_0_in1_data;
	wire cst_0_in1_ready;
	wire cst_0_in1_valid;
	wire [0 : 0]cst_0_out1_data;
	wire cst_0_out1_ready;
	wire cst_0_out1_valid;

	wire branch_0_clk;
	wire branch_0_rst;
	wire [0 : 0]branch_0_in1_data;
	wire branch_0_in1_ready;
	wire branch_0_in1_valid;
	wire [0 : 0]branch_0_in2_data;
	wire branch_0_in2_ready;
	wire branch_0_in2_valid;
	wire [0 : 0]branch_0_out1_data;
	wire branch_0_out1_ready;
	wire branch_0_out1_valid;
	wire [0 : 0]branch_0_out2_data;
	wire branch_0_out2_ready;
	wire branch_0_out2_valid;

	wire start_0_clk;
	wire start_0_rst;
	wire [0 : 0]start_0_in1_data;
	wire start_0_in1_ready;
	wire start_0_in1_valid;
	wire [0 : 0]start_0_out1_data;
	wire start_0_out1_ready;
	wire start_0_out1_valid;

	wire forkC_24_clk;
	wire forkC_24_rst;
	wire [0 : 0]forkC_24_in1_data;
	wire forkC_24_in1_ready;
	wire forkC_24_in1_valid;
	wire [0 : 0]forkC_24_out1_data;
	wire forkC_24_out1_ready;
	wire forkC_24_out1_valid;
	wire [0 : 0]forkC_24_out2_data;
	wire forkC_24_out2_ready;
	wire forkC_24_out2_valid;
	wire [0 : 0]forkC_24_out3_data;
	wire forkC_24_out3_ready;
	wire forkC_24_out3_valid;

	wire branchC_26_clk;
	wire branchC_26_rst;
	wire [0 : 0]branchC_26_in1_data;
	wire branchC_26_in1_ready;
	wire branchC_26_in1_valid;
	wire [0 : 0]branchC_26_in2_data;
	wire branchC_26_in2_ready;
	wire branchC_26_in2_valid;
	wire [0 : 0]branchC_26_out1_data;
	wire branchC_26_out1_ready;
	wire branchC_26_out1_valid;
	wire [0 : 0]branchC_26_out2_data;
	wire branchC_26_out2_ready;
	wire branchC_26_out2_valid;

	wire fork_25_clk;
	wire fork_25_rst;
	wire [0 : 0]fork_25_in1_data;
	wire fork_25_in1_ready;
	wire fork_25_in1_valid;
	wire [0 : 0]fork_25_out1_data;
	wire fork_25_out1_ready;
	wire fork_25_out1_valid;
	wire [0 : 0]fork_25_out2_data;
	wire fork_25_out2_ready;
	wire fork_25_out2_valid;

	wire MC_filter_clk;
	wire MC_filter_rst;
	wire [5 : 0]MC_filter_in1_data;
	wire MC_filter_in1_ready;
	wire MC_filter_in1_valid;
	wire [31 : 0]MC_filter_in2_data;
	wire MC_filter_in2_ready;
	wire MC_filter_in2_valid;
	wire [5 : 0]MC_filter_in3_data;
	wire MC_filter_in3_ready;
	wire MC_filter_in3_valid;
	wire [31 : 0]MC_filter_in4_data;
	wire MC_filter_in4_ready;
	wire MC_filter_in4_valid;
	wire [31 : 0]MC_filter_out1_data;
	wire MC_filter_out1_ready;
	wire MC_filter_out1_valid;
	wire [0 : 0]MC_filter_out2_data;
	wire MC_filter_out2_ready;
	wire MC_filter_out2_valid;

	wire MC_orig_clk;
	wire MC_orig_rst;
	wire [12 : 0]MC_orig_in1_data;
	wire MC_orig_in1_ready;
	wire MC_orig_in1_valid;
	wire [31 : 0]MC_orig_in2_data;
	wire MC_orig_in2_ready;
	wire MC_orig_in2_valid;
	wire [12 : 0]MC_orig_in3_data;
	wire MC_orig_in3_ready;
	wire MC_orig_in3_valid;
	wire [31 : 0]MC_orig_in4_data;
	wire MC_orig_in4_ready;
	wire MC_orig_in4_valid;
	wire [31 : 0]MC_orig_out1_data;
	wire MC_orig_out1_ready;
	wire MC_orig_out1_valid;
	wire [0 : 0]MC_orig_out2_data;
	wire MC_orig_out2_ready;
	wire MC_orig_out2_valid;

	wire MC_sol_clk;
	wire MC_sol_rst;
	wire [31 : 0]MC_sol_in1_data;
	wire MC_sol_in1_ready;
	wire MC_sol_in1_valid;
	wire [10 : 0]MC_sol_in2_data;
	wire MC_sol_in2_ready;
	wire MC_sol_in2_valid;
	wire [31 : 0]MC_sol_in3_data;
	wire MC_sol_in3_ready;
	wire MC_sol_in3_valid;
	wire [10 : 0]MC_sol_in4_data;
	wire MC_sol_in4_ready;
	wire MC_sol_in4_valid;
	wire [0 : 0]MC_sol_out1_data;
	wire MC_sol_out1_ready;
	wire MC_sol_out1_valid;
	wire [31 : 0]MC_sol_out2_data;
	wire MC_sol_out2_ready;
	wire MC_sol_out2_valid;

	wire sink_1_clk;
	wire sink_1_rst;
	wire [0 : 0]sink_1_in1_data;
	wire sink_1_in1_ready;
	wire sink_1_in1_valid;

	wire sink_2_clk;
	wire sink_2_rst;
	wire [0 : 0]sink_2_in1_data;
	wire sink_2_in1_ready;
	wire sink_2_in1_valid;

	wire sink_3_clk;
	wire sink_3_rst;
	wire [4 : 0]sink_3_in1_data;
	wire sink_3_in1_ready;
	wire sink_3_in1_valid;

	wire sink_4_clk;
	wire sink_4_rst;
	wire [0 : 0]sink_4_in1_data;
	wire sink_4_in1_ready;
	wire sink_4_in1_valid;

	wire sink_5_clk;
	wire sink_5_rst;
	wire [0 : 0]sink_5_in1_data;
	wire sink_5_in1_ready;
	wire sink_5_in1_valid;

	wire sink_6_clk;
	wire sink_6_rst;
	wire [4 : 0]sink_6_in1_data;
	wire sink_6_in1_ready;
	wire sink_6_in1_valid;

	wire sink_7_clk;
	wire sink_7_rst;
	wire [4 : 0]sink_7_in1_data;
	wire sink_7_in1_ready;
	wire sink_7_in1_valid;

	wire sink_8_clk;
	wire sink_8_rst;
	wire [0 : 0]sink_8_in1_data;
	wire sink_8_in1_ready;
	wire sink_8_in1_valid;

	wire sink_9_clk;
	wire sink_9_rst;
	wire [31 : 0]sink_9_in1_data;
	wire sink_9_in1_ready;
	wire sink_9_in1_valid;

	wire sink_10_clk;
	wire sink_10_rst;
	wire [2 : 0]sink_10_in1_data;
	wire sink_10_in1_ready;
	wire sink_10_in1_valid;

	wire sink_11_clk;
	wire sink_11_rst;
	wire [4 : 0]sink_11_in1_data;
	wire sink_11_in1_ready;
	wire sink_11_in1_valid;

	wire sink_12_clk;
	wire sink_12_rst;
	wire [4 : 0]sink_12_in1_data;
	wire sink_12_in1_ready;
	wire sink_12_in1_valid;

	wire sink_13_clk;
	wire sink_13_rst;
	wire [2 : 0]sink_13_in1_data;
	wire sink_13_in1_ready;
	wire sink_13_in1_valid;

	wire sink_14_clk;
	wire sink_14_rst;
	wire [2 : 0]sink_14_in1_data;
	wire sink_14_in1_ready;
	wire sink_14_in1_valid;

	wire sink_15_clk;
	wire sink_15_rst;
	wire [4 : 0]sink_15_in1_data;
	wire sink_15_in1_ready;
	wire sink_15_in1_valid;

	wire sink_16_clk;
	wire sink_16_rst;
	wire [31 : 0]sink_16_in1_data;
	wire sink_16_in1_ready;
	wire sink_16_in1_valid;

	wire sink_17_clk;
	wire sink_17_rst;
	wire [31 : 0]sink_17_in1_data;
	wire sink_17_in1_ready;
	wire sink_17_in1_valid;

	wire sink_18_clk;
	wire sink_18_rst;
	wire [4 : 0]sink_18_in1_data;
	wire sink_18_in1_ready;
	wire sink_18_in1_valid;

	wire sink_19_clk;
	wire sink_19_rst;
	wire [0 : 0]sink_19_in1_data;
	wire sink_19_in1_ready;
	wire sink_19_in1_valid;

	wire sink_20_clk;
	wire sink_20_rst;
	wire [0 : 0]sink_20_in1_data;
	wire sink_20_in1_ready;
	wire sink_20_in1_valid;

	wire sink_21_clk;
	wire sink_21_rst;
	wire [0 : 0]sink_21_in1_data;
	wire sink_21_in1_ready;
	wire sink_21_in1_valid;

	wire sink_22_clk;
	wire sink_22_rst;
	wire [0 : 0]sink_22_in1_data;
	wire sink_22_in1_ready;
	wire sink_22_in1_valid;

	wire Buffer_100_clk;
	wire Buffer_100_rst;
	wire [31 : 0]Buffer_100_in1_data;
	wire Buffer_100_in1_ready;
	wire Buffer_100_in1_valid;
	wire [31 : 0]Buffer_100_out1_data;
	wire Buffer_100_out1_ready;
	wire Buffer_100_out1_valid;

	wire Buffer_101_clk;
	wire Buffer_101_rst;
	wire [31 : 0]Buffer_101_in1_data;
	wire Buffer_101_in1_ready;
	wire Buffer_101_in1_valid;
	wire [31 : 0]Buffer_101_out1_data;
	wire Buffer_101_out1_ready;
	wire Buffer_101_out1_valid;

	wire Buffer_102_clk;
	wire Buffer_102_rst;
	wire [31 : 0]Buffer_102_in1_data;
	wire Buffer_102_in1_ready;
	wire Buffer_102_in1_valid;
	wire [31 : 0]Buffer_102_out1_data;
	wire Buffer_102_out1_ready;
	wire Buffer_102_out1_valid;

	wire Buffer_103_clk;
	wire Buffer_103_rst;
	wire [31 : 0]Buffer_103_in1_data;
	wire Buffer_103_in1_ready;
	wire Buffer_103_in1_valid;
	wire [31 : 0]Buffer_103_out1_data;
	wire Buffer_103_out1_ready;
	wire Buffer_103_out1_valid;

	wire Buffer_104_clk;
	wire Buffer_104_rst;
	wire [31 : 0]Buffer_104_in1_data;
	wire Buffer_104_in1_ready;
	wire Buffer_104_in1_valid;
	wire [31 : 0]Buffer_104_out1_data;
	wire Buffer_104_out1_ready;
	wire Buffer_104_out1_valid;

	wire Buffer_105_clk;
	wire Buffer_105_rst;
	wire [31 : 0]Buffer_105_in1_data;
	wire Buffer_105_in1_ready;
	wire Buffer_105_in1_valid;
	wire [31 : 0]Buffer_105_out1_data;
	wire Buffer_105_out1_ready;
	wire Buffer_105_out1_valid;

	wire Buffer_106_clk;
	wire Buffer_106_rst;
	wire [31 : 0]Buffer_106_in1_data;
	wire Buffer_106_in1_ready;
	wire Buffer_106_in1_valid;
	wire [31 : 0]Buffer_106_out1_data;
	wire Buffer_106_out1_ready;
	wire Buffer_106_out1_valid;

	wire Buffer_107_clk;
	wire Buffer_107_rst;
	wire [31 : 0]Buffer_107_in1_data;
	wire Buffer_107_in1_ready;
	wire Buffer_107_in1_valid;
	wire [31 : 0]Buffer_107_out1_data;
	wire Buffer_107_out1_ready;
	wire Buffer_107_out1_valid;

	wire Buffer_108_clk;
	wire Buffer_108_rst;
	wire [31 : 0]Buffer_108_in1_data;
	wire Buffer_108_in1_ready;
	wire Buffer_108_in1_valid;
	wire [31 : 0]Buffer_108_out1_data;
	wire Buffer_108_out1_ready;
	wire Buffer_108_out1_valid;

	wire Buffer_109_clk;
	wire Buffer_109_rst;
	wire [31 : 0]Buffer_109_in1_data;
	wire Buffer_109_in1_ready;
	wire Buffer_109_in1_valid;
	wire [31 : 0]Buffer_109_out1_data;
	wire Buffer_109_out1_ready;
	wire Buffer_109_out1_valid;

	wire Buffer_110_clk;
	wire Buffer_110_rst;
	wire [31 : 0]Buffer_110_in1_data;
	wire Buffer_110_in1_ready;
	wire Buffer_110_in1_valid;
	wire [31 : 0]Buffer_110_out1_data;
	wire Buffer_110_out1_ready;
	wire Buffer_110_out1_valid;

	wire Buffer_111_clk;
	wire Buffer_111_rst;
	wire [31 : 0]Buffer_111_in1_data;
	wire Buffer_111_in1_ready;
	wire Buffer_111_in1_valid;
	wire [31 : 0]Buffer_111_out1_data;
	wire Buffer_111_out1_ready;
	wire Buffer_111_out1_valid;

	wire Buffer_112_clk;
	wire Buffer_112_rst;
	wire [31 : 0]Buffer_112_in1_data;
	wire Buffer_112_in1_ready;
	wire Buffer_112_in1_valid;
	wire [31 : 0]Buffer_112_out1_data;
	wire Buffer_112_out1_ready;
	wire Buffer_112_out1_valid;

	wire Buffer_113_clk;
	wire Buffer_113_rst;
	wire [31 : 0]Buffer_113_in1_data;
	wire Buffer_113_in1_ready;
	wire Buffer_113_in1_valid;
	wire [31 : 0]Buffer_113_out1_data;
	wire Buffer_113_out1_ready;
	wire Buffer_113_out1_valid;

	wire Buffer_114_clk;
	wire Buffer_114_rst;
	wire [31 : 0]Buffer_114_in1_data;
	wire Buffer_114_in1_ready;
	wire Buffer_114_in1_valid;
	wire [31 : 0]Buffer_114_out1_data;
	wire Buffer_114_out1_ready;
	wire Buffer_114_out1_valid;

	wire Buffer_115_clk;
	wire Buffer_115_rst;
	wire [31 : 0]Buffer_115_in1_data;
	wire Buffer_115_in1_ready;
	wire Buffer_115_in1_valid;
	wire [31 : 0]Buffer_115_out1_data;
	wire Buffer_115_out1_ready;
	wire Buffer_115_out1_valid;



	assign phi_5_clk = clk;
	assign phi_5_rst = rst;
	assign branch_9_in1_data = phi_5_out1_data;
	assign branch_9_in1_valid = phi_5_out1_valid;
	assign phi_5_out1_ready = branch_9_in1_ready;

	assign phi_6_clk = clk;
	assign phi_6_rst = rst;
	assign branch_8_in1_data = phi_6_out1_data;
	assign branch_8_in1_valid = phi_6_out1_valid;
	assign phi_6_out1_ready = branch_8_in1_ready;

	assign brCst_block4_clk = clk;
	assign brCst_block4_rst = rst;
	assign fork_18_in1_data = brCst_block4_out1_data;
	assign fork_18_in1_valid = brCst_block4_out1_valid;
	assign brCst_block4_out1_ready = fork_18_in1_ready;

	assign cst_4_clk = clk;
	assign cst_4_rst = rst;
	assign branch_7_in1_data = cst_4_out1_data;
	assign branch_7_in1_valid = cst_4_out1_valid;
	assign cst_4_out1_ready = branch_7_in1_ready;

	assign phi_n6_clk = clk;
	assign phi_n6_rst = rst;
	assign branch_10_in1_data = phi_n6_out1_data;
	assign branch_10_in1_valid = phi_n6_out1_valid;
	assign phi_n6_out1_ready = branch_10_in1_ready;

	assign phi_n7_clk = clk;
	assign phi_n7_rst = rst;
	assign branch_11_in1_data = phi_n7_out1_data;
	assign branch_11_in1_valid = phi_n7_out1_valid;
	assign phi_n7_out1_ready = branch_11_in1_ready;

	assign branch_7_clk = clk;
	assign branch_7_rst = rst;
	assign phi_8_in2_data = branch_7_out1_data;
	assign phi_8_in2_valid = branch_7_out1_valid;
	assign branch_7_out1_ready = phi_8_in2_ready;
	assign sink_8_in1_data = branch_7_out2_data;
	assign sink_8_in1_valid = branch_7_out2_valid;
	assign branch_7_out2_ready = sink_8_in1_ready;

	assign branch_8_clk = clk;
	assign branch_8_rst = rst;
	assign phi_9_in2_data = branch_8_out1_data;
	assign phi_9_in2_valid = branch_8_out1_valid;
	assign branch_8_out1_ready = phi_9_in2_ready;
	assign sink_9_in1_data = branch_8_out2_data;
	assign sink_9_in1_valid = branch_8_out2_valid;
	assign branch_8_out2_ready = sink_9_in1_ready;

	assign branch_9_clk = clk;
	assign branch_9_rst = rst;
	assign phi_n12_in1_data = branch_9_out1_data;
	assign phi_n12_in1_valid = branch_9_out1_valid;
	assign branch_9_out1_ready = phi_n12_in1_ready;
	assign sink_10_in1_data = branch_9_out2_data;
	assign sink_10_in1_valid = branch_9_out2_valid;
	assign branch_9_out2_ready = sink_10_in1_ready;

	assign branch_10_clk = clk;
	assign branch_10_rst = rst;
	assign phi_n13_in1_data = branch_10_out1_data;
	assign phi_n13_in1_valid = branch_10_out1_valid;
	assign branch_10_out1_ready = phi_n13_in1_ready;
	assign sink_11_in1_data = branch_10_out2_data;
	assign sink_11_in1_valid = branch_10_out2_valid;
	assign branch_10_out2_ready = sink_11_in1_ready;

	assign branch_11_clk = clk;
	assign branch_11_rst = rst;
	assign phi_n14_in1_data = branch_11_out1_data;
	assign phi_n14_in1_valid = branch_11_out1_valid;
	assign branch_11_out1_ready = phi_n14_in1_ready;
	assign sink_12_in1_data = branch_11_out2_data;
	assign sink_12_in1_valid = branch_11_out2_valid;
	assign branch_11_out2_ready = sink_12_in1_ready;

	assign fork_18_clk = clk;
	assign fork_18_rst = rst;
	assign branch_11_in2_data = fork_18_out1_data;
	assign branch_11_in2_valid = fork_18_out1_valid;
	assign fork_18_out1_ready = branch_11_in2_ready;
	assign branch_10_in2_data = fork_18_out2_data;
	assign branch_10_in2_valid = fork_18_out2_valid;
	assign fork_18_out2_ready = branch_10_in2_ready;
	assign branch_9_in2_data = fork_18_out3_data;
	assign branch_9_in2_valid = fork_18_out3_valid;
	assign fork_18_out3_ready = branch_9_in2_ready;
	assign branch_8_in2_data = fork_18_out4_data;
	assign branch_8_in2_valid = fork_18_out4_valid;
	assign fork_18_out4_ready = branch_8_in2_ready;
	assign branch_7_in2_data = fork_18_out5_data;
	assign branch_7_in2_valid = fork_18_out5_valid;
	assign fork_18_out5_ready = branch_7_in2_ready;
	assign branchC_29_in2_data = fork_18_out6_data;
	assign branchC_29_in2_valid = fork_18_out6_valid;
	assign fork_18_out6_ready = branchC_29_in2_ready;

	assign phiC_18_clk = clk;
	assign phiC_18_rst = rst;
	assign forkC_28_in1_data = phiC_18_out1_data;
	assign forkC_28_in1_valid = phiC_18_out1_valid;
	assign phiC_18_out1_ready = forkC_28_in1_ready;
	assign fork_36_in1_data = phiC_18_out2_data;
	assign fork_36_in1_valid = phiC_18_out2_valid;
	assign phiC_18_out2_ready = fork_36_in1_ready;

	assign forkC_28_clk = clk;
	assign forkC_28_rst = rst;
	assign cst_4_in1_data = forkC_28_out1_data;
	assign cst_4_in1_valid = forkC_28_out1_valid;
	assign forkC_28_out1_ready = cst_4_in1_ready;
	assign branchC_29_in1_data = forkC_28_out2_data;
	assign branchC_29_in1_valid = forkC_28_out2_valid;
	assign forkC_28_out2_ready = branchC_29_in1_ready;
	assign brCst_block4_in1_data = forkC_28_out3_data;
	assign brCst_block4_in1_valid = forkC_28_out3_valid;
	assign forkC_28_out3_ready = brCst_block4_in1_ready;

	assign branchC_29_clk = clk;
	assign branchC_29_rst = rst;
	assign phiC_19_in1_data = branchC_29_out1_data;
	assign phiC_19_in1_valid = branchC_29_out1_valid;
	assign branchC_29_out1_ready = phiC_19_in1_ready;
	assign sink_22_in1_data = branchC_29_out2_data;
	assign sink_22_in1_valid = branchC_29_out2_valid;
	assign branchC_29_out2_ready = sink_22_in1_ready;

	assign fork_36_clk = clk;
	assign fork_36_rst = rst;
	assign phi_5_in1_data = fork_36_out1_data;
	assign phi_5_in1_valid = fork_36_out1_valid;
	assign fork_36_out1_ready = phi_5_in1_ready;
	assign phi_6_in1_data = fork_36_out2_data;
	assign phi_6_in1_valid = fork_36_out2_valid;
	assign fork_36_out2_ready = phi_6_in1_ready;

	assign cst_9_clk = clk;
	assign cst_9_rst = rst;
	assign add_27_in2_data = cst_9_out1_data;
	assign add_27_in2_valid = cst_9_out1_valid;
	assign cst_9_out1_ready = add_27_in2_ready;

	assign add_27_clk = clk;
	assign add_27_rst = rst;
	assign fork_3_in1_data = add_27_out1_data;
	assign fork_3_in1_valid = add_27_out1_valid;
	assign add_27_out1_ready = fork_3_in1_ready;

	assign cst_10_clk = clk;
	assign cst_10_rst = rst;
	assign icmp_28_in2_data = cst_10_out1_data;
	assign icmp_28_in2_valid = cst_10_out1_valid;
	assign cst_10_out1_ready = icmp_28_in2_ready;

	assign icmp_28_clk = clk;
	assign icmp_28_rst = rst;
	assign fork_20_in1_data = icmp_28_out1_data;
	assign fork_20_in1_valid = icmp_28_out1_valid;
	assign icmp_28_out1_ready = fork_20_in1_ready;

	assign phi_n8_clk = clk;
	assign phi_n8_rst = rst;
	assign add_27_in1_data = phi_n8_out1_data;
	assign add_27_in1_valid = phi_n8_out1_valid;
	assign phi_n8_out1_ready = add_27_in1_ready;

	assign phi_n9_clk = clk;
	assign phi_n9_rst = rst;
	assign branch_18_in1_data = phi_n9_out1_data;
	assign branch_18_in1_valid = phi_n9_out1_valid;
	assign phi_n9_out1_ready = branch_18_in1_ready;

	assign phi_n10_clk = clk;
	assign phi_n10_rst = rst;
	assign branch_19_in1_data = phi_n10_out1_data;
	assign branch_19_in1_valid = phi_n10_out1_valid;
	assign phi_n10_out1_ready = branch_19_in1_ready;

	assign phi_n11_clk = clk;
	assign phi_n11_rst = rst;
	assign branch_20_in1_data = phi_n11_out1_data;
	assign branch_20_in1_valid = phi_n11_out1_valid;
	assign phi_n11_out1_ready = branch_20_in1_ready;

	assign fork_3_clk = clk;
	assign fork_3_rst = rst;
	assign icmp_28_in1_data = fork_3_out1_data;
	assign icmp_28_in1_valid = fork_3_out1_valid;
	assign fork_3_out1_ready = icmp_28_in1_ready;
	assign branch_17_in1_data = fork_3_out2_data;
	assign branch_17_in1_valid = fork_3_out2_valid;
	assign fork_3_out2_ready = branch_17_in1_ready;

	assign branch_17_clk = clk;
	assign branch_17_rst = rst;
	assign Buffer_106_in1_data = branch_17_out1_data;
	assign Buffer_106_in1_valid = branch_17_out1_valid;
	assign branch_17_out1_ready = Buffer_106_in1_ready;
	assign sink_14_in1_data = branch_17_out2_data;
	assign sink_14_in1_valid = branch_17_out2_valid;
	assign branch_17_out2_ready = sink_14_in1_ready;

	assign branch_18_clk = clk;
	assign branch_18_rst = rst;
	assign Buffer_107_in1_data = branch_18_out1_data;
	assign Buffer_107_in1_valid = branch_18_out1_valid;
	assign branch_18_out1_ready = Buffer_107_in1_ready;
	assign phi_n5_in1_data = branch_18_out2_data;
	assign phi_n5_in1_valid = branch_18_out2_valid;
	assign branch_18_out2_ready = phi_n5_in1_ready;

	assign branch_19_clk = clk;
	assign branch_19_rst = rst;
	assign Buffer_108_in1_data = branch_19_out1_data;
	assign Buffer_108_in1_valid = branch_19_out1_valid;
	assign branch_19_out1_ready = Buffer_108_in1_ready;
	assign phi_n3_in1_data = branch_19_out2_data;
	assign phi_n3_in1_valid = branch_19_out2_valid;
	assign branch_19_out2_ready = phi_n3_in1_ready;

	assign branch_20_clk = clk;
	assign branch_20_rst = rst;
	assign Buffer_109_in1_data = branch_20_out1_data;
	assign Buffer_109_in1_valid = branch_20_out1_valid;
	assign branch_20_out1_ready = Buffer_109_in1_ready;
	assign phi_n4_in1_data = branch_20_out2_data;
	assign phi_n4_in1_valid = branch_20_out2_valid;
	assign branch_20_out2_ready = phi_n4_in1_ready;

	assign fork_20_clk = clk;
	assign fork_20_rst = rst;
	assign branch_20_in2_data = fork_20_out1_data;
	assign branch_20_in2_valid = fork_20_out1_valid;
	assign fork_20_out1_ready = branch_20_in2_ready;
	assign branch_19_in2_data = fork_20_out2_data;
	assign branch_19_in2_valid = fork_20_out2_valid;
	assign fork_20_out2_ready = branch_19_in2_ready;
	assign branch_18_in2_data = fork_20_out3_data;
	assign branch_18_in2_valid = fork_20_out3_valid;
	assign fork_20_out3_ready = branch_18_in2_ready;
	assign branch_17_in2_data = fork_20_out4_data;
	assign branch_17_in2_valid = fork_20_out4_valid;
	assign fork_20_out4_ready = branch_17_in2_ready;
	assign branchC_31_in2_data = fork_20_out5_data;
	assign branchC_31_in2_valid = fork_20_out5_valid;
	assign fork_20_out5_ready = branchC_31_in2_ready;

	assign phiC_20_clk = clk;
	assign phiC_20_rst = rst;
	assign branchC_31_in1_data = phiC_20_out1_data;
	assign branchC_31_in1_valid = phiC_20_out1_valid;
	assign phiC_20_out1_ready = branchC_31_in1_ready;

	assign branchC_31_clk = clk;
	assign branchC_31_rst = rst;
	assign Buffer_110_in1_data = branchC_31_out1_data;
	assign Buffer_110_in1_valid = branchC_31_out1_valid;
	assign branchC_31_out1_ready = Buffer_110_in1_ready;
	assign phiC_21_in1_data = branchC_31_out2_data;
	assign phiC_21_in1_valid = branchC_31_out2_valid;
	assign branchC_31_out2_ready = phiC_21_in1_ready;

	assign source_4_clk = clk;
	assign source_4_rst = rst;
	assign cst_9_in1_data = source_4_out1_data;
	assign cst_9_in1_valid = source_4_out1_valid;
	assign source_4_out1_ready = cst_9_in1_ready;

	assign source_5_clk = clk;
	assign source_5_rst = rst;
	assign cst_10_in1_data = source_5_out1_data;
	assign cst_10_in1_valid = source_5_out1_valid;
	assign source_5_out1_ready = cst_10_in1_ready;

	assign cst_14_clk = clk;
	assign cst_14_rst = rst;
	assign add_37_in2_data = cst_14_out1_data;
	assign add_37_in2_valid = cst_14_out1_valid;
	assign cst_14_out1_ready = add_37_in2_ready;

	assign add_37_clk = clk;
	assign add_37_rst = rst;
	assign fork_5_in1_data = add_37_out1_data;
	assign fork_5_in1_valid = add_37_out1_valid;
	assign add_37_out1_ready = fork_5_in1_ready;

	assign cst_15_clk = clk;
	assign cst_15_rst = rst;
	assign icmp_38_in2_data = cst_15_out1_data;
	assign icmp_38_in2_valid = cst_15_out1_valid;
	assign cst_15_out1_ready = icmp_38_in2_ready;

	assign icmp_38_clk = clk;
	assign icmp_38_rst = rst;
	assign fork_22_in1_data = icmp_38_out1_data;
	assign fork_22_in1_valid = icmp_38_out1_valid;
	assign icmp_38_out1_ready = fork_22_in1_ready;

	assign phi_n0_clk = clk;
	assign phi_n0_rst = rst;
	assign add_37_in1_data = phi_n0_out1_data;
	assign add_37_in1_valid = phi_n0_out1_valid;
	assign phi_n0_out1_ready = add_37_in1_ready;

	assign phi_n1_clk = clk;
	assign phi_n1_rst = rst;
	assign branch_24_in1_data = phi_n1_out1_data;
	assign branch_24_in1_valid = phi_n1_out1_valid;
	assign phi_n1_out1_ready = branch_24_in1_ready;

	assign fork_5_clk = clk;
	assign fork_5_rst = rst;
	assign icmp_38_in1_data = fork_5_out1_data;
	assign icmp_38_in1_valid = fork_5_out1_valid;
	assign fork_5_out1_ready = icmp_38_in1_ready;
	assign branch_25_in1_data = fork_5_out2_data;
	assign branch_25_in1_valid = fork_5_out2_valid;
	assign fork_5_out2_ready = branch_25_in1_ready;

	assign branch_24_clk = clk;
	assign branch_24_rst = rst;
	assign sink_17_in1_data = branch_24_out1_data;
	assign sink_17_in1_valid = branch_24_out1_valid;
	assign branch_24_out1_ready = sink_17_in1_ready;
	assign phi_n15_in1_data = branch_24_out2_data;
	assign phi_n15_in1_valid = branch_24_out2_valid;
	assign branch_24_out2_ready = phi_n15_in1_ready;

	assign branch_25_clk = clk;
	assign branch_25_rst = rst;
	assign Buffer_114_in1_data = branch_25_out1_data;
	assign Buffer_114_in1_valid = branch_25_out1_valid;
	assign branch_25_out1_ready = Buffer_114_in1_ready;
	assign sink_18_in1_data = branch_25_out2_data;
	assign sink_18_in1_valid = branch_25_out2_valid;
	assign branch_25_out2_ready = sink_18_in1_ready;

	assign fork_22_clk = clk;
	assign fork_22_rst = rst;
	assign branch_25_in2_data = fork_22_out1_data;
	assign branch_25_in2_valid = fork_22_out1_valid;
	assign fork_22_out1_ready = branch_25_in2_ready;
	assign branch_24_in2_data = fork_22_out2_data;
	assign branch_24_in2_valid = fork_22_out2_valid;
	assign fork_22_out2_ready = branch_24_in2_ready;
	assign branchC_33_in2_data = fork_22_out3_data;
	assign branchC_33_in2_valid = fork_22_out3_valid;
	assign fork_22_out3_ready = branchC_33_in2_ready;

	assign phiC_22_clk = clk;
	assign phiC_22_rst = rst;
	assign branchC_33_in1_data = phiC_22_out1_data;
	assign branchC_33_in1_valid = phiC_22_out1_valid;
	assign phiC_22_out1_ready = branchC_33_in1_ready;

	assign branchC_33_clk = clk;
	assign branchC_33_rst = rst;
	assign Buffer_115_in1_data = branchC_33_out1_data;
	assign Buffer_115_in1_valid = branchC_33_out1_valid;
	assign branchC_33_out1_ready = Buffer_115_in1_ready;
	assign phiC_23_in1_data = branchC_33_out2_data;
	assign phiC_23_in1_valid = branchC_33_out2_valid;
	assign branchC_33_out2_ready = phiC_23_in1_ready;

	assign source_9_clk = clk;
	assign source_9_rst = rst;
	assign cst_14_in1_data = source_9_out1_data;
	assign cst_14_in1_valid = source_9_out1_valid;
	assign source_9_out1_ready = cst_14_in1_ready;

	assign source_10_clk = clk;
	assign source_10_rst = rst;
	assign cst_15_in1_data = source_10_out1_data;
	assign cst_15_in1_valid = source_10_out1_valid;
	assign source_10_out1_ready = cst_15_in1_ready;

	assign ret_0_clk = clk;
	assign ret_0_rst = rst;
	assign end_0_in4_data = ret_0_out1_data;
	assign end_0_in4_valid = ret_0_out1_valid;
	assign ret_0_out1_ready = end_0_in4_ready;

	assign phi_n15_clk = clk;
	assign phi_n15_rst = rst;
	assign ret_0_in1_data = phi_n15_out1_data;
	assign ret_0_in1_valid = phi_n15_out1_valid;
	assign phi_n15_out1_ready = ret_0_in1_ready;

	assign end_0_clk = clk;
	assign end_0_rst = rst;
	assign end_out = end_0_out1_data;
	assign end_0_out1_ready = end_ready;
	assign end_valid = end_0_out1_valid;

	assign phiC_23_clk = clk;
	assign phiC_23_rst = rst;
	assign sink_0_in1_data = phiC_23_out1_data;
	assign sink_0_in1_valid = phiC_23_out1_valid;
	assign phiC_23_out1_ready = sink_0_in1_ready;

	assign sink_0_clk = clk;
	assign sink_0_rst = rst;

	assign phi_3_clk = clk;
	assign phi_3_rst = rst;
	assign branch_5_in1_data = phi_3_out1_data;
	assign branch_5_in1_valid = phi_3_out1_valid;
	assign phi_3_out1_ready = branch_5_in1_ready;

	assign brCst_block3_clk = clk;
	assign brCst_block3_rst = rst;
	assign fork_17_in1_data = brCst_block3_out1_data;
	assign fork_17_in1_valid = brCst_block3_out1_valid;
	assign brCst_block3_out1_ready = fork_17_in1_ready;

	assign cst_2_clk = clk;
	assign cst_2_rst = rst;
	assign branch_3_in1_data = cst_2_out1_data;
	assign branch_3_in1_valid = cst_2_out1_valid;
	assign cst_2_out1_ready = branch_3_in1_ready;

	assign cst_3_clk = clk;
	assign cst_3_rst = rst;
	assign branch_4_in1_data = cst_3_out1_data;
	assign branch_4_in1_valid = cst_3_out1_valid;
	assign cst_3_out1_ready = branch_4_in1_ready;

	assign phi_n2_clk = clk;
	assign phi_n2_rst = rst;
	assign branch_6_in1_data = phi_n2_out1_data;
	assign branch_6_in1_valid = phi_n2_out1_valid;
	assign phi_n2_out1_ready = branch_6_in1_ready;

	assign branch_3_clk = clk;
	assign branch_3_rst = rst;
	assign phi_5_in2_data = branch_3_out1_data;
	assign phi_5_in2_valid = branch_3_out1_valid;
	assign branch_3_out1_ready = phi_5_in2_ready;
	assign sink_4_in1_data = branch_3_out2_data;
	assign sink_4_in1_valid = branch_3_out2_valid;
	assign branch_3_out2_ready = sink_4_in1_ready;

	assign branch_4_clk = clk;
	assign branch_4_rst = rst;
	assign phi_6_in2_data = branch_4_out1_data;
	assign phi_6_in2_valid = branch_4_out1_valid;
	assign branch_4_out1_ready = phi_6_in2_ready;
	assign sink_5_in1_data = branch_4_out2_data;
	assign sink_5_in1_valid = branch_4_out2_valid;
	assign branch_4_out2_ready = sink_5_in1_ready;

	assign branch_5_clk = clk;
	assign branch_5_rst = rst;
	assign phi_n7_in1_data = branch_5_out1_data;
	assign phi_n7_in1_valid = branch_5_out1_valid;
	assign branch_5_out1_ready = phi_n7_in1_ready;
	assign sink_6_in1_data = branch_5_out2_data;
	assign sink_6_in1_valid = branch_5_out2_valid;
	assign branch_5_out2_ready = sink_6_in1_ready;

	assign branch_6_clk = clk;
	assign branch_6_rst = rst;
	assign phi_n6_in1_data = branch_6_out1_data;
	assign phi_n6_in1_valid = branch_6_out1_valid;
	assign branch_6_out1_ready = phi_n6_in1_ready;
	assign sink_7_in1_data = branch_6_out2_data;
	assign sink_7_in1_valid = branch_6_out2_valid;
	assign branch_6_out2_ready = sink_7_in1_ready;

	assign fork_17_clk = clk;
	assign fork_17_rst = rst;
	assign branch_6_in2_data = fork_17_out1_data;
	assign branch_6_in2_valid = fork_17_out1_valid;
	assign fork_17_out1_ready = branch_6_in2_ready;
	assign branch_5_in2_data = fork_17_out2_data;
	assign branch_5_in2_valid = fork_17_out2_valid;
	assign fork_17_out2_ready = branch_5_in2_ready;
	assign branch_4_in2_data = fork_17_out3_data;
	assign branch_4_in2_valid = fork_17_out3_valid;
	assign fork_17_out3_ready = branch_4_in2_ready;
	assign branch_3_in2_data = fork_17_out4_data;
	assign branch_3_in2_valid = fork_17_out4_valid;
	assign fork_17_out4_ready = branch_3_in2_ready;
	assign branchC_28_in2_data = fork_17_out5_data;
	assign branchC_28_in2_valid = fork_17_out5_valid;
	assign fork_17_out5_ready = branchC_28_in2_ready;

	assign phiC_17_clk = clk;
	assign phiC_17_rst = rst;
	assign forkC_27_in1_data = phiC_17_out1_data;
	assign forkC_27_in1_valid = phiC_17_out1_valid;
	assign phiC_17_out1_ready = forkC_27_in1_ready;
	assign phi_3_in1_data = phiC_17_out2_data;
	assign phi_3_in1_valid = phiC_17_out2_valid;
	assign phiC_17_out2_ready = phi_3_in1_ready;

	assign forkC_27_clk = clk;
	assign forkC_27_rst = rst;
	assign cst_2_in1_data = forkC_27_out1_data;
	assign cst_2_in1_valid = forkC_27_out1_valid;
	assign forkC_27_out1_ready = cst_2_in1_ready;
	assign cst_3_in1_data = forkC_27_out2_data;
	assign cst_3_in1_valid = forkC_27_out2_valid;
	assign forkC_27_out2_ready = cst_3_in1_ready;
	assign branchC_28_in1_data = forkC_27_out3_data;
	assign branchC_28_in1_valid = forkC_27_out3_valid;
	assign forkC_27_out3_ready = branchC_28_in1_ready;
	assign brCst_block3_in1_data = forkC_27_out4_data;
	assign brCst_block3_in1_valid = forkC_27_out4_valid;
	assign forkC_27_out4_ready = brCst_block3_in1_ready;

	assign branchC_28_clk = clk;
	assign branchC_28_rst = rst;
	assign phiC_18_in1_data = branchC_28_out1_data;
	assign phiC_18_in1_valid = branchC_28_out1_valid;
	assign branchC_28_out1_ready = phiC_18_in1_ready;
	assign sink_21_in1_data = branchC_28_out2_data;
	assign sink_21_in1_valid = branchC_28_out2_valid;
	assign branchC_28_out2_ready = sink_21_in1_ready;

	assign cst_11_clk = clk;
	assign cst_11_rst = rst;
	assign mul_30_in2_data = cst_11_out1_data;
	assign mul_30_in2_valid = cst_11_out1_valid;
	assign cst_11_out1_ready = mul_30_in2_ready;

	assign mul_30_clk = clk;
	assign mul_30_rst = rst;
	assign add_31_in1_data = mul_30_out1_data;
	assign add_31_in1_valid = mul_30_out1_valid;
	assign mul_30_out1_ready = add_31_in1_ready;

	assign add_31_clk = clk;
	assign add_31_rst = rst;
	assign store_0_in2_data = add_31_out1_data;
	assign store_0_in2_valid = add_31_out1_valid;
	assign add_31_out1_ready = store_0_in2_ready;

	assign store_0_clk = clk;
	assign store_0_rst = rst;
	assign MC_sol_in3_data = store_0_out1_data;
	assign MC_sol_in3_valid = store_0_out1_valid;
	assign store_0_out1_ready = MC_sol_in3_ready;
	assign MC_sol_in2_data = store_0_out2_data;
	assign MC_sol_in2_valid = store_0_out2_valid;
	assign store_0_out2_ready = MC_sol_in2_ready;

	assign cst_12_clk = clk;
	assign cst_12_rst = rst;
	assign add_34_in2_data = cst_12_out1_data;
	assign add_34_in2_valid = cst_12_out1_valid;
	assign cst_12_out1_ready = add_34_in2_ready;

	assign add_34_clk = clk;
	assign add_34_rst = rst;
	assign fork_4_in1_data = add_34_out1_data;
	assign fork_4_in1_valid = add_34_out1_valid;
	assign add_34_out1_ready = fork_4_in1_ready;

	assign cst_13_clk = clk;
	assign cst_13_rst = rst;
	assign icmp_35_in2_data = cst_13_out1_data;
	assign icmp_35_in2_valid = cst_13_out1_valid;
	assign cst_13_out1_ready = icmp_35_in2_ready;

	assign icmp_35_clk = clk;
	assign icmp_35_rst = rst;
	assign fork_21_in1_data = icmp_35_out1_data;
	assign fork_21_in1_valid = icmp_35_out1_valid;
	assign icmp_35_out1_ready = fork_21_in1_ready;

	assign phi_n3_clk = clk;
	assign phi_n3_rst = rst;
	assign fork_6_in1_data = phi_n3_out1_data;
	assign fork_6_in1_valid = phi_n3_out1_valid;
	assign phi_n3_out1_ready = fork_6_in1_ready;

	assign phi_n4_clk = clk;
	assign phi_n4_rst = rst;
	assign fork_7_in1_data = phi_n4_out1_data;
	assign fork_7_in1_valid = phi_n4_out1_valid;
	assign phi_n4_out1_ready = fork_7_in1_ready;

	assign phi_n5_clk = clk;
	assign phi_n5_rst = rst;
	assign fork_8_in1_data = phi_n5_out1_data;
	assign fork_8_in1_valid = phi_n5_out1_valid;
	assign phi_n5_out1_ready = fork_8_in1_ready;

	assign fork_4_clk = clk;
	assign fork_4_rst = rst;
	assign icmp_35_in1_data = fork_4_out1_data;
	assign icmp_35_in1_valid = fork_4_out1_valid;
	assign fork_4_out1_ready = icmp_35_in1_ready;
	assign branch_21_in1_data = fork_4_out2_data;
	assign branch_21_in1_valid = fork_4_out2_valid;
	assign fork_4_out2_ready = branch_21_in1_ready;

	assign fork_6_clk = clk;
	assign fork_6_rst = rst;
	assign mul_30_in1_data = fork_6_out1_data;
	assign mul_30_in1_valid = fork_6_out1_valid;
	assign fork_6_out1_ready = mul_30_in1_ready;
	assign branch_22_in1_data = fork_6_out2_data;
	assign branch_22_in1_valid = fork_6_out2_valid;
	assign fork_6_out2_ready = branch_22_in1_ready;

	assign fork_7_clk = clk;
	assign fork_7_rst = rst;
	assign add_31_in2_data = fork_7_out1_data;
	assign add_31_in2_valid = fork_7_out1_valid;
	assign fork_7_out1_ready = add_31_in2_ready;
	assign add_34_in1_data = fork_7_out2_data;
	assign add_34_in1_valid = fork_7_out2_valid;
	assign fork_7_out2_ready = add_34_in1_ready;

	assign fork_8_clk = clk;
	assign fork_8_rst = rst;
	assign store_0_in1_data = fork_8_out1_data;
	assign store_0_in1_valid = fork_8_out1_valid;
	assign fork_8_out1_ready = store_0_in1_ready;
	assign branch_23_in1_data = fork_8_out2_data;
	assign branch_23_in1_valid = fork_8_out2_valid;
	assign fork_8_out2_ready = branch_23_in1_ready;

	assign branch_21_clk = clk;
	assign branch_21_rst = rst;
	assign Buffer_111_in1_data = branch_21_out1_data;
	assign Buffer_111_in1_valid = branch_21_out1_valid;
	assign branch_21_out1_ready = Buffer_111_in1_ready;
	assign sink_15_in1_data = branch_21_out2_data;
	assign sink_15_in1_valid = branch_21_out2_valid;
	assign branch_21_out2_ready = sink_15_in1_ready;

	assign branch_22_clk = clk;
	assign branch_22_rst = rst;
	assign Buffer_112_in1_data = branch_22_out1_data;
	assign Buffer_112_in1_valid = branch_22_out1_valid;
	assign branch_22_out1_ready = Buffer_112_in1_ready;
	assign phi_n0_in1_data = branch_22_out2_data;
	assign phi_n0_in1_valid = branch_22_out2_valid;
	assign branch_22_out2_ready = phi_n0_in1_ready;

	assign branch_23_clk = clk;
	assign branch_23_rst = rst;
	assign sink_16_in1_data = branch_23_out1_data;
	assign sink_16_in1_valid = branch_23_out1_valid;
	assign branch_23_out1_ready = sink_16_in1_ready;
	assign phi_n1_in1_data = branch_23_out2_data;
	assign phi_n1_in1_valid = branch_23_out2_valid;
	assign branch_23_out2_ready = phi_n1_in1_ready;

	assign fork_21_clk = clk;
	assign fork_21_rst = rst;
	assign branch_23_in2_data = fork_21_out1_data;
	assign branch_23_in2_valid = fork_21_out1_valid;
	assign fork_21_out1_ready = branch_23_in2_ready;
	assign branch_22_in2_data = fork_21_out2_data;
	assign branch_22_in2_valid = fork_21_out2_valid;
	assign fork_21_out2_ready = branch_22_in2_ready;
	assign branch_21_in2_data = fork_21_out3_data;
	assign branch_21_in2_valid = fork_21_out3_valid;
	assign fork_21_out3_ready = branch_21_in2_ready;
	assign branchC_32_in2_data = fork_21_out4_data;
	assign branchC_32_in2_valid = fork_21_out4_valid;
	assign fork_21_out4_ready = branchC_32_in2_ready;

	assign cst_16_clk = clk;
	assign cst_16_rst = rst;
	assign MC_sol_in1_data = cst_16_out1_data;
	assign MC_sol_in1_valid = cst_16_out1_valid;
	assign cst_16_out1_ready = MC_sol_in1_ready;

	assign phiC_21_clk = clk;
	assign phiC_21_rst = rst;
	assign forkC_31_in1_data = phiC_21_out1_data;
	assign forkC_31_in1_valid = phiC_21_out1_valid;
	assign phiC_21_out1_ready = forkC_31_in1_ready;

	assign forkC_31_clk = clk;
	assign forkC_31_rst = rst;
	assign cst_16_in1_data = forkC_31_out1_data;
	assign cst_16_in1_valid = forkC_31_out1_valid;
	assign forkC_31_out1_ready = cst_16_in1_ready;
	assign branchC_32_in1_data = forkC_31_out2_data;
	assign branchC_32_in1_valid = forkC_31_out2_valid;
	assign forkC_31_out2_ready = branchC_32_in1_ready;

	assign branchC_32_clk = clk;
	assign branchC_32_rst = rst;
	assign Buffer_113_in1_data = branchC_32_out1_data;
	assign Buffer_113_in1_valid = branchC_32_out1_valid;
	assign branchC_32_out1_ready = Buffer_113_in1_ready;
	assign phiC_22_in1_data = branchC_32_out2_data;
	assign phiC_22_in1_valid = branchC_32_out2_valid;
	assign branchC_32_out2_ready = phiC_22_in1_ready;

	assign source_6_clk = clk;
	assign source_6_rst = rst;
	assign cst_11_in1_data = source_6_out1_data;
	assign cst_11_in1_valid = source_6_out1_valid;
	assign source_6_out1_ready = cst_11_in1_ready;

	assign source_7_clk = clk;
	assign source_7_rst = rst;
	assign cst_12_in1_data = source_7_out1_data;
	assign cst_12_in1_valid = source_7_out1_valid;
	assign source_7_out1_ready = cst_12_in1_ready;

	assign source_8_clk = clk;
	assign source_8_rst = rst;
	assign cst_13_in1_data = source_8_out1_data;
	assign cst_13_in1_valid = source_8_out1_valid;
	assign source_8_out1_ready = cst_13_in1_ready;

	assign phi_1_clk = clk;
	assign phi_1_rst = rst;
	assign branch_2_in1_data = phi_1_out1_data;
	assign branch_2_in1_valid = phi_1_out1_valid;
	assign phi_1_out1_ready = branch_2_in1_ready;

	assign brCst_block2_clk = clk;
	assign brCst_block2_rst = rst;
	assign fork_16_in1_data = brCst_block2_out1_data;
	assign fork_16_in1_valid = brCst_block2_out1_valid;
	assign brCst_block2_out1_ready = fork_16_in1_ready;

	assign cst_1_clk = clk;
	assign cst_1_rst = rst;
	assign branch_1_in1_data = cst_1_out1_data;
	assign branch_1_in1_valid = cst_1_out1_valid;
	assign cst_1_out1_ready = branch_1_in1_ready;

	assign branch_1_clk = clk;
	assign branch_1_rst = rst;
	assign phi_3_in2_data = branch_1_out1_data;
	assign phi_3_in2_valid = branch_1_out1_valid;
	assign branch_1_out1_ready = phi_3_in2_ready;
	assign sink_2_in1_data = branch_1_out2_data;
	assign sink_2_in1_valid = branch_1_out2_valid;
	assign branch_1_out2_ready = sink_2_in1_ready;

	assign branch_2_clk = clk;
	assign branch_2_rst = rst;
	assign phi_n2_in1_data = branch_2_out1_data;
	assign phi_n2_in1_valid = branch_2_out1_valid;
	assign branch_2_out1_ready = phi_n2_in1_ready;
	assign sink_3_in1_data = branch_2_out2_data;
	assign sink_3_in1_valid = branch_2_out2_valid;
	assign branch_2_out2_ready = sink_3_in1_ready;

	assign fork_16_clk = clk;
	assign fork_16_rst = rst;
	assign branch_2_in2_data = fork_16_out1_data;
	assign branch_2_in2_valid = fork_16_out1_valid;
	assign fork_16_out1_ready = branch_2_in2_ready;
	assign branch_1_in2_data = fork_16_out2_data;
	assign branch_1_in2_valid = fork_16_out2_valid;
	assign fork_16_out2_ready = branch_1_in2_ready;
	assign branchC_27_in2_data = fork_16_out3_data;
	assign branchC_27_in2_valid = fork_16_out3_valid;
	assign fork_16_out3_ready = branchC_27_in2_ready;

	assign phiC_16_clk = clk;
	assign phiC_16_rst = rst;
	assign forkC_26_in1_data = phiC_16_out1_data;
	assign forkC_26_in1_valid = phiC_16_out1_valid;
	assign phiC_16_out1_ready = forkC_26_in1_ready;
	assign phi_1_in1_data = phiC_16_out2_data;
	assign phi_1_in1_valid = phiC_16_out2_valid;
	assign phiC_16_out2_ready = phi_1_in1_ready;

	assign forkC_26_clk = clk;
	assign forkC_26_rst = rst;
	assign cst_1_in1_data = forkC_26_out1_data;
	assign cst_1_in1_valid = forkC_26_out1_valid;
	assign forkC_26_out1_ready = cst_1_in1_ready;
	assign branchC_27_in1_data = forkC_26_out2_data;
	assign branchC_27_in1_valid = forkC_26_out2_valid;
	assign forkC_26_out2_ready = branchC_27_in1_ready;
	assign brCst_block2_in1_data = forkC_26_out3_data;
	assign brCst_block2_in1_valid = forkC_26_out3_valid;
	assign forkC_26_out3_ready = brCst_block2_in1_ready;

	assign branchC_27_clk = clk;
	assign branchC_27_rst = rst;
	assign phiC_17_in1_data = branchC_27_out1_data;
	assign phiC_17_in1_valid = branchC_27_out1_valid;
	assign branchC_27_out1_ready = phiC_17_in1_ready;
	assign sink_20_in1_data = branchC_27_out2_data;
	assign sink_20_in1_valid = branchC_27_out2_valid;
	assign branchC_27_out2_ready = sink_20_in1_ready;

	assign phi_8_clk = clk;
	assign phi_8_rst = rst;
	assign fork_0_in1_data = phi_8_out1_data;
	assign fork_0_in1_valid = phi_8_out1_valid;
	assign phi_8_out1_ready = fork_0_in1_ready;

	assign phi_9_clk = clk;
	assign phi_9_rst = rst;
	assign add_23_in1_data = phi_9_out1_data;
	assign add_23_in1_valid = phi_9_out1_valid;
	assign phi_9_out1_ready = add_23_in1_ready;

	assign cst_5_clk = clk;
	assign cst_5_rst = rst;
	assign mul_10_in2_data = cst_5_out1_data;
	assign mul_10_in2_valid = cst_5_out1_valid;
	assign cst_5_out1_ready = mul_10_in2_ready;

	assign mul_10_clk = clk;
	assign mul_10_rst = rst;
	assign add_11_in1_data = mul_10_out1_data;
	assign add_11_in1_valid = mul_10_out1_valid;
	assign mul_10_out1_ready = add_11_in1_ready;

	assign add_11_clk = clk;
	assign add_11_rst = rst;
	assign load_14_in2_data = add_11_out1_data;
	assign load_14_in2_valid = add_11_out1_valid;
	assign add_11_out1_ready = load_14_in2_ready;

	assign load_14_clk = clk;
	assign load_14_rst = rst;
	assign mul_22_in1_data = load_14_out1_data;
	assign mul_22_in1_valid = load_14_out1_valid;
	assign load_14_out1_ready = mul_22_in1_ready;
	assign MC_filter_in1_data = load_14_out2_data;
	assign MC_filter_in1_valid = load_14_out2_valid;
	assign load_14_out2_ready = MC_filter_in1_ready;

	assign add_15_clk = clk;
	assign add_15_rst = rst;
	assign mul_16_in1_data = add_15_out1_data;
	assign mul_16_in1_valid = add_15_out1_valid;
	assign add_15_out1_ready = mul_16_in1_ready;

	assign cst_6_clk = clk;
	assign cst_6_rst = rst;
	assign mul_16_in2_data = cst_6_out1_data;
	assign mul_16_in2_valid = cst_6_out1_valid;
	assign cst_6_out1_ready = mul_16_in2_ready;

	assign mul_16_clk = clk;
	assign mul_16_rst = rst;
	assign add_17_in1_data = mul_16_out1_data;
	assign add_17_in1_valid = mul_16_out1_valid;
	assign mul_16_out1_ready = add_17_in1_ready;

	assign add_17_clk = clk;
	assign add_17_rst = rst;
	assign add_18_in1_data = add_17_out1_data;
	assign add_18_in1_valid = add_17_out1_valid;
	assign add_17_out1_ready = add_18_in1_ready;

	assign add_18_clk = clk;
	assign add_18_rst = rst;
	assign load_21_in2_data = add_18_out1_data;
	assign load_21_in2_valid = add_18_out1_valid;
	assign add_18_out1_ready = load_21_in2_ready;

	assign load_21_clk = clk;
	assign load_21_rst = rst;
	assign mul_22_in2_data = load_21_out1_data;
	assign mul_22_in2_valid = load_21_out1_valid;
	assign load_21_out1_ready = mul_22_in2_ready;
	assign MC_orig_in1_data = load_21_out2_data;
	assign MC_orig_in1_valid = load_21_out2_valid;
	assign load_21_out2_ready = MC_orig_in1_ready;

	assign mul_22_clk = clk;
	assign mul_22_rst = rst;
	assign add_23_in2_data = mul_22_out1_data;
	assign add_23_in2_valid = mul_22_out1_valid;
	assign mul_22_out1_ready = add_23_in2_ready;

	assign add_23_clk = clk;
	assign add_23_rst = rst;
	assign branch_12_in1_data = add_23_out1_data;
	assign branch_12_in1_valid = add_23_out1_valid;
	assign add_23_out1_ready = branch_12_in1_ready;

	assign cst_7_clk = clk;
	assign cst_7_rst = rst;
	assign add_24_in2_data = cst_7_out1_data;
	assign add_24_in2_valid = cst_7_out1_valid;
	assign cst_7_out1_ready = add_24_in2_ready;

	assign add_24_clk = clk;
	assign add_24_rst = rst;
	assign fork_2_in1_data = add_24_out1_data;
	assign fork_2_in1_valid = add_24_out1_valid;
	assign add_24_out1_ready = fork_2_in1_ready;

	assign cst_8_clk = clk;
	assign cst_8_rst = rst;
	assign icmp_25_in2_data = cst_8_out1_data;
	assign icmp_25_in2_valid = cst_8_out1_valid;
	assign cst_8_out1_ready = icmp_25_in2_ready;

	assign icmp_25_clk = clk;
	assign icmp_25_rst = rst;
	assign fork_19_in1_data = icmp_25_out1_data;
	assign fork_19_in1_valid = icmp_25_out1_valid;
	assign icmp_25_out1_ready = fork_19_in1_ready;

	assign phi_n12_clk = clk;
	assign phi_n12_rst = rst;
	assign fork_12_in1_data = phi_n12_out1_data;
	assign fork_12_in1_valid = phi_n12_out1_valid;
	assign phi_n12_out1_ready = fork_12_in1_ready;

	assign phi_n13_clk = clk;
	assign phi_n13_rst = rst;
	assign fork_13_in1_data = phi_n13_out1_data;
	assign fork_13_in1_valid = phi_n13_out1_valid;
	assign phi_n13_out1_ready = fork_13_in1_ready;

	assign phi_n14_clk = clk;
	assign phi_n14_rst = rst;
	assign fork_14_in1_data = phi_n14_out1_data;
	assign fork_14_in1_valid = phi_n14_out1_valid;
	assign phi_n14_out1_ready = fork_14_in1_ready;

	assign fork_0_clk = clk;
	assign fork_0_rst = rst;
	assign add_11_in2_data = fork_0_out1_data;
	assign add_11_in2_valid = fork_0_out1_valid;
	assign fork_0_out1_ready = add_11_in2_ready;
	assign add_18_in2_data = fork_0_out2_data;
	assign add_18_in2_valid = fork_0_out2_valid;
	assign fork_0_out2_ready = add_18_in2_ready;
	assign add_24_in1_data = fork_0_out3_data;
	assign add_24_in1_valid = fork_0_out3_valid;
	assign fork_0_out3_ready = add_24_in1_ready;

	assign fork_2_clk = clk;
	assign fork_2_rst = rst;
	assign icmp_25_in1_data = fork_2_out1_data;
	assign icmp_25_in1_valid = fork_2_out1_valid;
	assign fork_2_out1_ready = icmp_25_in1_ready;
	assign branch_13_in1_data = fork_2_out2_data;
	assign branch_13_in1_valid = fork_2_out2_valid;
	assign fork_2_out2_ready = branch_13_in1_ready;

	assign fork_12_clk = clk;
	assign fork_12_rst = rst;
	assign mul_10_in1_data = fork_12_out1_data;
	assign mul_10_in1_valid = fork_12_out1_valid;
	assign fork_12_out1_ready = mul_10_in1_ready;
	assign add_15_in2_data = fork_12_out2_data;
	assign add_15_in2_valid = fork_12_out2_valid;
	assign fork_12_out2_ready = add_15_in2_ready;
	assign branch_14_in1_data = fork_12_out3_data;
	assign branch_14_in1_valid = fork_12_out3_valid;
	assign fork_12_out3_ready = branch_14_in1_ready;

	assign fork_13_clk = clk;
	assign fork_13_rst = rst;
	assign add_15_in1_data = fork_13_out1_data;
	assign add_15_in1_valid = fork_13_out1_valid;
	assign fork_13_out1_ready = add_15_in1_ready;
	assign branch_15_in1_data = fork_13_out2_data;
	assign branch_15_in1_valid = fork_13_out2_valid;
	assign fork_13_out2_ready = branch_15_in1_ready;

	assign fork_14_clk = clk;
	assign fork_14_rst = rst;
	assign add_17_in2_data = fork_14_out1_data;
	assign add_17_in2_valid = fork_14_out1_valid;
	assign fork_14_out1_ready = add_17_in2_ready;
	assign branch_16_in1_data = fork_14_out2_data;
	assign branch_16_in1_valid = fork_14_out2_valid;
	assign fork_14_out2_ready = branch_16_in1_ready;

	assign branch_12_clk = clk;
	assign branch_12_rst = rst;
	assign Buffer_100_in1_data = branch_12_out1_data;
	assign Buffer_100_in1_valid = branch_12_out1_valid;
	assign branch_12_out1_ready = Buffer_100_in1_ready;
	assign phi_n9_in1_data = branch_12_out2_data;
	assign phi_n9_in1_valid = branch_12_out2_valid;
	assign branch_12_out2_ready = phi_n9_in1_ready;

	assign branch_13_clk = clk;
	assign branch_13_rst = rst;
	assign Buffer_101_in1_data = branch_13_out1_data;
	assign Buffer_101_in1_valid = branch_13_out1_valid;
	assign branch_13_out1_ready = Buffer_101_in1_ready;
	assign sink_13_in1_data = branch_13_out2_data;
	assign sink_13_in1_valid = branch_13_out2_valid;
	assign branch_13_out2_ready = sink_13_in1_ready;

	assign branch_14_clk = clk;
	assign branch_14_rst = rst;
	assign Buffer_102_in1_data = branch_14_out1_data;
	assign Buffer_102_in1_valid = branch_14_out1_valid;
	assign branch_14_out1_ready = Buffer_102_in1_ready;
	assign phi_n8_in1_data = branch_14_out2_data;
	assign phi_n8_in1_valid = branch_14_out2_valid;
	assign branch_14_out2_ready = phi_n8_in1_ready;

	assign branch_15_clk = clk;
	assign branch_15_rst = rst;
	assign Buffer_103_in1_data = branch_15_out1_data;
	assign Buffer_103_in1_valid = branch_15_out1_valid;
	assign branch_15_out1_ready = Buffer_103_in1_ready;
	assign phi_n10_in1_data = branch_15_out2_data;
	assign phi_n10_in1_valid = branch_15_out2_valid;
	assign branch_15_out2_ready = phi_n10_in1_ready;

	assign branch_16_clk = clk;
	assign branch_16_rst = rst;
	assign Buffer_104_in1_data = branch_16_out1_data;
	assign Buffer_104_in1_valid = branch_16_out1_valid;
	assign branch_16_out1_ready = Buffer_104_in1_ready;
	assign phi_n11_in1_data = branch_16_out2_data;
	assign phi_n11_in1_valid = branch_16_out2_valid;
	assign branch_16_out2_ready = phi_n11_in1_ready;

	assign fork_19_clk = clk;
	assign fork_19_rst = rst;
	assign branch_16_in2_data = fork_19_out1_data;
	assign branch_16_in2_valid = fork_19_out1_valid;
	assign fork_19_out1_ready = branch_16_in2_ready;
	assign branch_15_in2_data = fork_19_out2_data;
	assign branch_15_in2_valid = fork_19_out2_valid;
	assign fork_19_out2_ready = branch_15_in2_ready;
	assign branch_14_in2_data = fork_19_out3_data;
	assign branch_14_in2_valid = fork_19_out3_valid;
	assign fork_19_out3_ready = branch_14_in2_ready;
	assign branch_13_in2_data = fork_19_out4_data;
	assign branch_13_in2_valid = fork_19_out4_valid;
	assign fork_19_out4_ready = branch_13_in2_ready;
	assign branch_12_in2_data = fork_19_out5_data;
	assign branch_12_in2_valid = fork_19_out5_valid;
	assign fork_19_out5_ready = branch_12_in2_ready;
	assign branchC_30_in2_data = fork_19_out6_data;
	assign branchC_30_in2_valid = fork_19_out6_valid;
	assign fork_19_out6_ready = branchC_30_in2_ready;

	assign phiC_19_clk = clk;
	assign phiC_19_rst = rst;
	assign branchC_30_in1_data = phiC_19_out1_data;
	assign branchC_30_in1_valid = phiC_19_out1_valid;
	assign phiC_19_out1_ready = branchC_30_in1_ready;
	assign fork_37_in1_data = phiC_19_out2_data;
	assign fork_37_in1_valid = phiC_19_out2_valid;
	assign phiC_19_out2_ready = fork_37_in1_ready;

	assign branchC_30_clk = clk;
	assign branchC_30_rst = rst;
	assign Buffer_105_in1_data = branchC_30_out1_data;
	assign Buffer_105_in1_valid = branchC_30_out1_valid;
	assign branchC_30_out1_ready = Buffer_105_in1_ready;
	assign phiC_20_in1_data = branchC_30_out2_data;
	assign phiC_20_in1_valid = branchC_30_out2_valid;
	assign branchC_30_out2_ready = phiC_20_in1_ready;

	assign source_0_clk = clk;
	assign source_0_rst = rst;
	assign cst_5_in1_data = source_0_out1_data;
	assign cst_5_in1_valid = source_0_out1_valid;
	assign source_0_out1_ready = cst_5_in1_ready;

	assign source_1_clk = clk;
	assign source_1_rst = rst;
	assign cst_6_in1_data = source_1_out1_data;
	assign cst_6_in1_valid = source_1_out1_valid;
	assign source_1_out1_ready = cst_6_in1_ready;

	assign source_2_clk = clk;
	assign source_2_rst = rst;
	assign cst_7_in1_data = source_2_out1_data;
	assign cst_7_in1_valid = source_2_out1_valid;
	assign source_2_out1_ready = cst_7_in1_ready;

	assign source_3_clk = clk;
	assign source_3_rst = rst;
	assign cst_8_in1_data = source_3_out1_data;
	assign cst_8_in1_valid = source_3_out1_valid;
	assign source_3_out1_ready = cst_8_in1_ready;

	assign fork_37_clk = clk;
	assign fork_37_rst = rst;
	assign phi_8_in1_data = fork_37_out1_data;
	assign phi_8_in1_valid = fork_37_out1_valid;
	assign fork_37_out1_ready = phi_8_in1_ready;
	assign phi_9_in1_data = fork_37_out2_data;
	assign phi_9_in1_valid = fork_37_out2_valid;
	assign fork_37_out2_ready = phi_9_in1_ready;

	assign brCst_block1_clk = clk;
	assign brCst_block1_rst = rst;
	assign fork_25_in1_data = brCst_block1_out1_data;
	assign fork_25_in1_valid = brCst_block1_out1_valid;
	assign brCst_block1_out1_ready = fork_25_in1_ready;

	assign cst_0_clk = clk;
	assign cst_0_rst = rst;
	assign branch_0_in1_data = cst_0_out1_data;
	assign branch_0_in1_valid = cst_0_out1_valid;
	assign cst_0_out1_ready = branch_0_in1_ready;

	assign branch_0_clk = clk;
	assign branch_0_rst = rst;
	assign phi_1_in2_data = branch_0_out1_data;
	assign phi_1_in2_valid = branch_0_out1_valid;
	assign branch_0_out1_ready = phi_1_in2_ready;
	assign sink_1_in1_data = branch_0_out2_data;
	assign sink_1_in1_valid = branch_0_out2_valid;
	assign branch_0_out2_ready = sink_1_in1_ready;

	assign start_0_clk = clk;
	assign start_0_rst = rst;
	assign start_0_in1_data = start_in;
	assign start_0_in1_valid = start_valid;
	assign start_ready = start_0_in1_ready;
	assign forkC_24_in1_data = start_0_out1_data;
	assign forkC_24_in1_valid = start_0_out1_valid;
	assign start_0_out1_ready = forkC_24_in1_ready;

	assign forkC_24_clk = clk;
	assign forkC_24_rst = rst;
	assign cst_0_in1_data = forkC_24_out1_data;
	assign cst_0_in1_valid = forkC_24_out1_valid;
	assign forkC_24_out1_ready = cst_0_in1_ready;
	assign branchC_26_in1_data = forkC_24_out2_data;
	assign branchC_26_in1_valid = forkC_24_out2_valid;
	assign forkC_24_out2_ready = branchC_26_in1_ready;
	assign brCst_block1_in1_data = forkC_24_out3_data;
	assign brCst_block1_in1_valid = forkC_24_out3_valid;
	assign forkC_24_out3_ready = brCst_block1_in1_ready;

	assign branchC_26_clk = clk;
	assign branchC_26_rst = rst;
	assign phiC_16_in1_data = branchC_26_out1_data;
	assign phiC_16_in1_valid = branchC_26_out1_valid;
	assign branchC_26_out1_ready = phiC_16_in1_ready;
	assign sink_19_in1_data = branchC_26_out2_data;
	assign sink_19_in1_valid = branchC_26_out2_valid;
	assign branchC_26_out2_ready = sink_19_in1_ready;

	assign fork_25_clk = clk;
	assign fork_25_rst = rst;
	assign branch_0_in2_data = fork_25_out1_data;
	assign branch_0_in2_valid = fork_25_out1_valid;
	assign fork_25_out1_ready = branch_0_in2_ready;
	assign branchC_26_in2_data = fork_25_out2_data;
	assign branchC_26_in2_valid = fork_25_out2_valid;
	assign fork_25_out2_ready = branchC_26_in2_ready;

	assign MC_filter_clk = clk;
	assign MC_filter_rst = rst;
	assign filter_ce0 = filter_we0;
	assign MC_filter_in2_valid = 0;
	assign MC_filter_in2_data = 0;
	assign load_14_in1_data = MC_filter_out1_data;
	assign load_14_in1_valid = MC_filter_out1_valid;
	assign MC_filter_out1_ready = load_14_in1_ready;
	assign end_0_in1_data = MC_filter_out2_data;
	assign end_0_in1_valid = MC_filter_out2_valid;
	assign MC_filter_out2_ready = end_0_in1_ready;

	assign MC_orig_clk = clk;
	assign MC_orig_rst = rst;
	assign orig_ce0 = orig_we0;
	assign MC_orig_in2_valid = 0;
	assign MC_orig_in2_data = 0;
	assign load_21_in1_data = MC_orig_out1_data;
	assign load_21_in1_valid = MC_orig_out1_valid;
	assign MC_orig_out1_ready = load_21_in1_ready;
	assign end_0_in2_data = MC_orig_out2_data;
	assign end_0_in2_valid = MC_orig_out2_valid;
	assign MC_orig_out2_ready = end_0_in2_ready;

	assign MC_sol_clk = clk;
	assign MC_sol_rst = rst;
	assign sol_ce0 = sol_we0;
	assign end_0_in3_data = MC_sol_out1_data;
	assign end_0_in3_valid = MC_sol_out1_valid;
	assign MC_sol_out1_ready = end_0_in3_ready;

	assign sink_1_clk = clk;
	assign sink_1_rst = rst;

	assign sink_2_clk = clk;
	assign sink_2_rst = rst;

	assign sink_3_clk = clk;
	assign sink_3_rst = rst;

	assign sink_4_clk = clk;
	assign sink_4_rst = rst;

	assign sink_5_clk = clk;
	assign sink_5_rst = rst;

	assign sink_6_clk = clk;
	assign sink_6_rst = rst;

	assign sink_7_clk = clk;
	assign sink_7_rst = rst;

	assign sink_8_clk = clk;
	assign sink_8_rst = rst;

	assign sink_9_clk = clk;
	assign sink_9_rst = rst;

	assign sink_10_clk = clk;
	assign sink_10_rst = rst;

	assign sink_11_clk = clk;
	assign sink_11_rst = rst;

	assign sink_12_clk = clk;
	assign sink_12_rst = rst;

	assign sink_13_clk = clk;
	assign sink_13_rst = rst;

	assign sink_14_clk = clk;
	assign sink_14_rst = rst;

	assign sink_15_clk = clk;
	assign sink_15_rst = rst;

	assign sink_16_clk = clk;
	assign sink_16_rst = rst;

	assign sink_17_clk = clk;
	assign sink_17_rst = rst;

	assign sink_18_clk = clk;
	assign sink_18_rst = rst;

	assign sink_19_clk = clk;
	assign sink_19_rst = rst;

	assign sink_20_clk = clk;
	assign sink_20_rst = rst;

	assign sink_21_clk = clk;
	assign sink_21_rst = rst;

	assign sink_22_clk = clk;
	assign sink_22_rst = rst;

	assign Buffer_100_clk = clk;
	assign Buffer_100_rst = rst;
	assign phi_9_in3_data = Buffer_100_out1_data;
	assign phi_9_in3_valid = Buffer_100_out1_valid;
	assign Buffer_100_out1_ready = phi_9_in3_ready;

	assign Buffer_101_clk = clk;
	assign Buffer_101_rst = rst;
	assign phi_8_in3_data = Buffer_101_out1_data;
	assign phi_8_in3_valid = Buffer_101_out1_valid;
	assign Buffer_101_out1_ready = phi_8_in3_ready;

	assign Buffer_102_clk = clk;
	assign Buffer_102_rst = rst;
	assign phi_n12_in2_data = Buffer_102_out1_data;
	assign phi_n12_in2_valid = Buffer_102_out1_valid;
	assign Buffer_102_out1_ready = phi_n12_in2_ready;

	assign Buffer_103_clk = clk;
	assign Buffer_103_rst = rst;
	assign phi_n13_in2_data = Buffer_103_out1_data;
	assign phi_n13_in2_valid = Buffer_103_out1_valid;
	assign Buffer_103_out1_ready = phi_n13_in2_ready;

	assign Buffer_104_clk = clk;
	assign Buffer_104_rst = rst;
	assign phi_n14_in2_data = Buffer_104_out1_data;
	assign phi_n14_in2_valid = Buffer_104_out1_valid;
	assign Buffer_104_out1_ready = phi_n14_in2_ready;

	assign Buffer_105_clk = clk;
	assign Buffer_105_rst = rst;
	assign phiC_19_in2_data = Buffer_105_out1_data;
	assign phiC_19_in2_valid = Buffer_105_out1_valid;
	assign Buffer_105_out1_ready = phiC_19_in2_ready;

	assign Buffer_106_clk = clk;
	assign Buffer_106_rst = rst;
	assign phi_5_in3_data = Buffer_106_out1_data;
	assign phi_5_in3_valid = Buffer_106_out1_valid;
	assign Buffer_106_out1_ready = phi_5_in3_ready;

	assign Buffer_107_clk = clk;
	assign Buffer_107_rst = rst;
	assign phi_6_in3_data = Buffer_107_out1_data;
	assign phi_6_in3_valid = Buffer_107_out1_valid;
	assign Buffer_107_out1_ready = phi_6_in3_ready;

	assign Buffer_108_clk = clk;
	assign Buffer_108_rst = rst;
	assign phi_n6_in2_data = Buffer_108_out1_data;
	assign phi_n6_in2_valid = Buffer_108_out1_valid;
	assign Buffer_108_out1_ready = phi_n6_in2_ready;

	assign Buffer_109_clk = clk;
	assign Buffer_109_rst = rst;
	assign phi_n7_in2_data = Buffer_109_out1_data;
	assign phi_n7_in2_valid = Buffer_109_out1_valid;
	assign Buffer_109_out1_ready = phi_n7_in2_ready;

	assign Buffer_110_clk = clk;
	assign Buffer_110_rst = rst;
	assign phiC_18_in2_data = Buffer_110_out1_data;
	assign phiC_18_in2_valid = Buffer_110_out1_valid;
	assign Buffer_110_out1_ready = phiC_18_in2_ready;

	assign Buffer_111_clk = clk;
	assign Buffer_111_rst = rst;
	assign phi_3_in3_data = Buffer_111_out1_data;
	assign phi_3_in3_valid = Buffer_111_out1_valid;
	assign Buffer_111_out1_ready = phi_3_in3_ready;

	assign Buffer_112_clk = clk;
	assign Buffer_112_rst = rst;
	assign phi_n2_in2_data = Buffer_112_out1_data;
	assign phi_n2_in2_valid = Buffer_112_out1_valid;
	assign Buffer_112_out1_ready = phi_n2_in2_ready;

	assign Buffer_113_clk = clk;
	assign Buffer_113_rst = rst;
	assign phiC_17_in2_data = Buffer_113_out1_data;
	assign phiC_17_in2_valid = Buffer_113_out1_valid;
	assign Buffer_113_out1_ready = phiC_17_in2_ready;

	assign Buffer_114_clk = clk;
	assign Buffer_114_rst = rst;
	assign phi_1_in3_data = Buffer_114_out1_data;
	assign phi_1_in3_valid = Buffer_114_out1_valid;
	assign Buffer_114_out1_ready = phi_1_in3_ready;

	assign Buffer_115_clk = clk;
	assign Buffer_115_rst = rst;
	assign phiC_16_in2_data = Buffer_115_out1_data;
	assign phiC_16_in2_valid = Buffer_115_out1_valid;
	assign Buffer_115_out1_ready = phiC_16_in2_ready;

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3), .COND_SIZE(1)) mux_node_phi_5
		(.clk(phi_5_clk), .rst(phi_5_rst),
		.data_in_bus({{2'b0, phi_5_in1_data}, phi_5_in3_data, phi_5_in2_data}), .valid_in_bus({phi_5_in1_valid, phi_5_in3_valid, phi_5_in2_valid}), .ready_in_bus({phi_5_in1_ready, phi_5_in3_ready, phi_5_in2_ready}), 
		.data_out_bus({phi_5_out1_data}), .valid_out_bus({phi_5_out1_valid}), .ready_out_bus({phi_5_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_6
		(.clk(phi_6_clk), .rst(phi_6_rst),
		.data_in_bus({{31'b0, phi_6_in1_data}, phi_6_in3_data, phi_6_in2_data}), .valid_in_bus({phi_6_in1_valid, phi_6_in3_valid, phi_6_in2_valid}), .ready_in_bus({phi_6_in1_ready, phi_6_in3_ready, phi_6_in2_ready}), 
		.data_out_bus({phi_6_out1_data}), .valid_out_bus({phi_6_out1_valid}), .ready_out_bus({phi_6_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block4
		(.clk(brCst_block4_clk), .rst(brCst_block4_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block4_in1_valid}), .ready_in_bus({brCst_block4_in1_ready}), 
		.data_out_bus({brCst_block4_out1_data}), .valid_out_bus({brCst_block4_out1_valid}), .ready_out_bus({brCst_block4_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_4
		(.clk(cst_4_clk), .rst(cst_4_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_4_in1_valid}), .ready_in_bus({cst_4_in1_ready}), 
		.data_out_bus({cst_4_out1_data}), .valid_out_bus({cst_4_out1_valid}), .ready_out_bus({cst_4_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n6
		(.clk(phi_n6_clk), .rst(phi_n6_rst),
		.data_in_bus({phi_n6_in2_data, phi_n6_in1_data}), .valid_in_bus({phi_n6_in2_valid, phi_n6_in1_valid}), .ready_in_bus({phi_n6_in2_ready, phi_n6_in1_ready}), 
		.data_out_bus({phi_n6_out1_data}), .valid_out_bus({phi_n6_out1_valid}), .ready_out_bus({phi_n6_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n7
		(.clk(phi_n7_clk), .rst(phi_n7_rst),
		.data_in_bus({phi_n7_in2_data, phi_n7_in1_data}), .valid_in_bus({phi_n7_in2_valid, phi_n7_in1_valid}), .ready_in_bus({phi_n7_in2_ready, phi_n7_in1_ready}), 
		.data_out_bus({phi_n7_out1_data}), .valid_out_bus({phi_n7_out1_valid}), .ready_out_bus({phi_n7_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_7
		(.clk(branch_7_clk), .rst(branch_7_rst),
		.data_in_bus({{branch_7_in2_data}, branch_7_in1_data}), .valid_in_bus({branch_7_in2_valid, branch_7_in1_valid}), .ready_in_bus({branch_7_in2_ready, branch_7_in1_ready}), 
		.data_out_bus({branch_7_out2_data, branch_7_out1_data}), .valid_out_bus({branch_7_out2_valid, branch_7_out1_valid}), .ready_out_bus({branch_7_out2_ready, branch_7_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_8
		(.clk(branch_8_clk), .rst(branch_8_rst),
		.data_in_bus({{31'b0, branch_8_in2_data}, branch_8_in1_data}), .valid_in_bus({branch_8_in2_valid, branch_8_in1_valid}), .ready_in_bus({branch_8_in2_ready, branch_8_in1_ready}), 
		.data_out_bus({branch_8_out2_data, branch_8_out1_data}), .valid_out_bus({branch_8_out2_valid, branch_8_out1_valid}), .ready_out_bus({branch_8_out2_ready, branch_8_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) branch_node_branch_9
		(.clk(branch_9_clk), .rst(branch_9_rst),
		.data_in_bus({{2'b0, branch_9_in2_data}, branch_9_in1_data}), .valid_in_bus({branch_9_in2_valid, branch_9_in1_valid}), .ready_in_bus({branch_9_in2_ready, branch_9_in1_ready}), 
		.data_out_bus({branch_9_out2_data, branch_9_out1_data}), .valid_out_bus({branch_9_out2_valid, branch_9_out1_valid}), .ready_out_bus({branch_9_out2_ready, branch_9_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_10
		(.clk(branch_10_clk), .rst(branch_10_rst),
		.data_in_bus({{4'b0, branch_10_in2_data}, branch_10_in1_data}), .valid_in_bus({branch_10_in2_valid, branch_10_in1_valid}), .ready_in_bus({branch_10_in2_ready, branch_10_in1_ready}), 
		.data_out_bus({branch_10_out2_data, branch_10_out1_data}), .valid_out_bus({branch_10_out2_valid, branch_10_out1_valid}), .ready_out_bus({branch_10_out2_ready, branch_10_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_11
		(.clk(branch_11_clk), .rst(branch_11_rst),
		.data_in_bus({{4'b0, branch_11_in2_data}, branch_11_in1_data}), .valid_in_bus({branch_11_in2_valid, branch_11_in1_valid}), .ready_in_bus({branch_11_in2_ready, branch_11_in1_ready}), 
		.data_out_bus({branch_11_out2_data, branch_11_out1_data}), .valid_out_bus({branch_11_out2_valid, branch_11_out1_valid}), .ready_out_bus({branch_11_out2_ready, branch_11_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(6), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_18
		(.clk(fork_18_clk), .rst(fork_18_rst),
		.data_in_bus({fork_18_in1_data}), .valid_in_bus({fork_18_in1_valid}), .ready_in_bus({fork_18_in1_ready}), 
		.data_out_bus({fork_18_out6_data, fork_18_out5_data, fork_18_out4_data, fork_18_out3_data, fork_18_out2_data, fork_18_out1_data}), .valid_out_bus({fork_18_out6_valid, fork_18_out5_valid, fork_18_out4_valid, fork_18_out3_valid, fork_18_out2_valid, fork_18_out1_valid}), .ready_out_bus({fork_18_out6_ready, fork_18_out5_ready, fork_18_out4_ready, fork_18_out3_ready, fork_18_out2_ready, fork_18_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_18
		(.clk(phiC_18_clk), .rst(phiC_18_rst),
		.data_in_bus({phiC_18_in2_data, phiC_18_in1_data}), .valid_in_bus({phiC_18_in2_valid, phiC_18_in1_valid}), .ready_in_bus({phiC_18_in2_ready, phiC_18_in1_ready}), 
		.data_out_bus({phiC_18_out2_data, phiC_18_out1_data}), .valid_out_bus({phiC_18_out2_valid, phiC_18_out1_valid}), .ready_out_bus({phiC_18_out2_ready, phiC_18_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_28
		(.clk(forkC_28_clk), .rst(forkC_28_rst),
		.data_in_bus({forkC_28_in1_data}), .valid_in_bus({forkC_28_in1_valid}), .ready_in_bus({forkC_28_in1_ready}), 
		.data_out_bus({forkC_28_out3_data, forkC_28_out2_data, forkC_28_out1_data}), .valid_out_bus({forkC_28_out3_valid, forkC_28_out2_valid, forkC_28_out1_valid}), .ready_out_bus({forkC_28_out3_ready, forkC_28_out2_ready, forkC_28_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_29
		(.clk(branchC_29_clk), .rst(branchC_29_rst),
		.data_in_bus({{branchC_29_in2_data}, branchC_29_in1_data}), .valid_in_bus({branchC_29_in2_valid, branchC_29_in1_valid}), .ready_in_bus({branchC_29_in2_ready, branchC_29_in1_ready}), 
		.data_out_bus({branchC_29_out2_data, branchC_29_out1_data}), .valid_out_bus({branchC_29_out2_valid, branchC_29_out1_valid}), .ready_out_bus({branchC_29_out2_ready, branchC_29_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_36
		(.clk(fork_36_clk), .rst(fork_36_rst),
		.data_in_bus({fork_36_in1_data}), .valid_in_bus({fork_36_in1_valid}), .ready_in_bus({fork_36_in1_ready}), 
		.data_out_bus({fork_36_out2_data, fork_36_out1_data}), .valid_out_bus({fork_36_out2_valid, fork_36_out1_valid}), .ready_out_bus({fork_36_out2_ready, fork_36_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_9
		(.clk(cst_9_clk), .rst(cst_9_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_9_in1_valid}), .ready_in_bus({cst_9_in1_ready}), 
		.data_out_bus({cst_9_out1_data}), .valid_out_bus({cst_9_out1_valid}), .ready_out_bus({cst_9_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) add_op_add_27
		(.clk(add_27_clk), .rst(add_27_rst),
		.data_in_bus({add_27_in2_data, add_27_in1_data}), .valid_in_bus({add_27_in2_valid, add_27_in1_valid}), .ready_in_bus({add_27_in2_ready, add_27_in1_ready}), 
		.data_out_bus({add_27_out1_data}), .valid_out_bus({add_27_out1_valid}), .ready_out_bus({add_27_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_10
		(.clk(cst_10_clk), .rst(cst_10_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_10_in1_valid}), .ready_in_bus({cst_10_in1_ready}), 
		.data_out_bus({cst_10_out1_data}), .valid_out_bus({cst_10_out1_valid}), .ready_out_bus({cst_10_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_28
		(.clk(icmp_28_clk), .rst(icmp_28_rst),
		.data_in_bus({icmp_28_in2_data, icmp_28_in1_data}), .valid_in_bus({icmp_28_in2_valid, icmp_28_in1_valid}), .ready_in_bus({icmp_28_in2_ready, icmp_28_in1_ready}), 
		.data_out_bus({icmp_28_out1_data}), .valid_out_bus({icmp_28_out1_valid}), .ready_out_bus({icmp_28_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) merge_node_phi_n8
		(.clk(phi_n8_clk), .rst(phi_n8_rst),
		.data_in_bus({phi_n8_in1_data}), .valid_in_bus({phi_n8_in1_valid}), .ready_in_bus({phi_n8_in1_ready}), 
		.data_out_bus({phi_n8_out1_data}), .valid_out_bus({phi_n8_out1_valid}), .ready_out_bus({phi_n8_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n9
		(.clk(phi_n9_clk), .rst(phi_n9_rst),
		.data_in_bus({phi_n9_in1_data}), .valid_in_bus({phi_n9_in1_valid}), .ready_in_bus({phi_n9_in1_ready}), 
		.data_out_bus({phi_n9_out1_data}), .valid_out_bus({phi_n9_out1_valid}), .ready_out_bus({phi_n9_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n10
		(.clk(phi_n10_clk), .rst(phi_n10_rst),
		.data_in_bus({phi_n10_in1_data}), .valid_in_bus({phi_n10_in1_valid}), .ready_in_bus({phi_n10_in1_ready}), 
		.data_out_bus({phi_n10_out1_data}), .valid_out_bus({phi_n10_out1_valid}), .ready_out_bus({phi_n10_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n11
		(.clk(phi_n11_clk), .rst(phi_n11_rst),
		.data_in_bus({phi_n11_in1_data}), .valid_in_bus({phi_n11_in1_valid}), .ready_in_bus({phi_n11_in1_ready}), 
		.data_out_bus({phi_n11_out1_data}), .valid_out_bus({phi_n11_out1_valid}), .ready_out_bus({phi_n11_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) fork_node_fork_3
		(.clk(fork_3_clk), .rst(fork_3_rst),
		.data_in_bus({fork_3_in1_data}), .valid_in_bus({fork_3_in1_valid}), .ready_in_bus({fork_3_in1_ready}), 
		.data_out_bus({fork_3_out2_data, fork_3_out1_data}), .valid_out_bus({fork_3_out2_valid, fork_3_out1_valid}), .ready_out_bus({fork_3_out2_ready, fork_3_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) branch_node_branch_17
		(.clk(branch_17_clk), .rst(branch_17_rst),
		.data_in_bus({{2'b0, branch_17_in2_data}, branch_17_in1_data}), .valid_in_bus({branch_17_in2_valid, branch_17_in1_valid}), .ready_in_bus({branch_17_in2_ready, branch_17_in1_ready}), 
		.data_out_bus({branch_17_out2_data, branch_17_out1_data}), .valid_out_bus({branch_17_out2_valid, branch_17_out1_valid}), .ready_out_bus({branch_17_out2_ready, branch_17_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_18
		(.clk(branch_18_clk), .rst(branch_18_rst),
		.data_in_bus({{31'b0, branch_18_in2_data}, branch_18_in1_data}), .valid_in_bus({branch_18_in2_valid, branch_18_in1_valid}), .ready_in_bus({branch_18_in2_ready, branch_18_in1_ready}), 
		.data_out_bus({branch_18_out2_data, branch_18_out1_data}), .valid_out_bus({branch_18_out2_valid, branch_18_out1_valid}), .ready_out_bus({branch_18_out2_ready, branch_18_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_19
		(.clk(branch_19_clk), .rst(branch_19_rst),
		.data_in_bus({{4'b0, branch_19_in2_data}, branch_19_in1_data}), .valid_in_bus({branch_19_in2_valid, branch_19_in1_valid}), .ready_in_bus({branch_19_in2_ready, branch_19_in1_ready}), 
		.data_out_bus({branch_19_out2_data, branch_19_out1_data}), .valid_out_bus({branch_19_out2_valid, branch_19_out1_valid}), .ready_out_bus({branch_19_out2_ready, branch_19_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_20
		(.clk(branch_20_clk), .rst(branch_20_rst),
		.data_in_bus({{4'b0, branch_20_in2_data}, branch_20_in1_data}), .valid_in_bus({branch_20_in2_valid, branch_20_in1_valid}), .ready_in_bus({branch_20_in2_ready, branch_20_in1_ready}), 
		.data_out_bus({branch_20_out2_data, branch_20_out1_data}), .valid_out_bus({branch_20_out2_valid, branch_20_out1_valid}), .ready_out_bus({branch_20_out2_ready, branch_20_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_20
		(.clk(fork_20_clk), .rst(fork_20_rst),
		.data_in_bus({fork_20_in1_data}), .valid_in_bus({fork_20_in1_valid}), .ready_in_bus({fork_20_in1_ready}), 
		.data_out_bus({fork_20_out5_data, fork_20_out4_data, fork_20_out3_data, fork_20_out2_data, fork_20_out1_data}), .valid_out_bus({fork_20_out5_valid, fork_20_out4_valid, fork_20_out3_valid, fork_20_out2_valid, fork_20_out1_valid}), .ready_out_bus({fork_20_out5_ready, fork_20_out4_ready, fork_20_out3_ready, fork_20_out2_ready, fork_20_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_20
		(.clk(phiC_20_clk), .rst(phiC_20_rst),
		.data_in_bus({phiC_20_in1_data}), .valid_in_bus({phiC_20_in1_valid}), .ready_in_bus({phiC_20_in1_ready}), 
		.data_out_bus({phiC_20_out1_data}), .valid_out_bus({phiC_20_out1_valid}), .ready_out_bus({phiC_20_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_31
		(.clk(branchC_31_clk), .rst(branchC_31_rst),
		.data_in_bus({{branchC_31_in2_data}, branchC_31_in1_data}), .valid_in_bus({branchC_31_in2_valid, branchC_31_in1_valid}), .ready_in_bus({branchC_31_in2_ready, branchC_31_in1_ready}), 
		.data_out_bus({branchC_31_out2_data, branchC_31_out1_data}), .valid_out_bus({branchC_31_out2_valid, branchC_31_out1_valid}), .ready_out_bus({branchC_31_out2_ready, branchC_31_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_4
		(.clk(source_4_clk), .rst(source_4_rst),
		.data_out_bus({source_4_out1_data}), .valid_out_bus({source_4_out1_valid}), .ready_out_bus({source_4_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_5
		(.clk(source_5_clk), .rst(source_5_rst),
		.data_out_bus({source_5_out1_data}), .valid_out_bus({source_5_out1_valid}), .ready_out_bus({source_5_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_14
		(.clk(cst_14_clk), .rst(cst_14_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_14_in1_valid}), .ready_in_bus({cst_14_in1_ready}), 
		.data_out_bus({cst_14_out1_data}), .valid_out_bus({cst_14_out1_valid}), .ready_out_bus({cst_14_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) add_op_add_37
		(.clk(add_37_clk), .rst(add_37_rst),
		.data_in_bus({add_37_in2_data, add_37_in1_data}), .valid_in_bus({add_37_in2_valid, add_37_in1_valid}), .ready_in_bus({add_37_in2_ready, add_37_in1_ready}), 
		.data_out_bus({add_37_out1_data}), .valid_out_bus({add_37_out1_valid}), .ready_out_bus({add_37_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) const_node_cst_15
		(.clk(cst_15_clk), .rst(cst_15_rst),
		.data_in_bus({5'd28}), .valid_in_bus({cst_15_in1_valid}), .ready_in_bus({cst_15_in1_ready}), 
		.data_out_bus({cst_15_out1_data}), .valid_out_bus({cst_15_out1_valid}), .ready_out_bus({cst_15_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_38
		(.clk(icmp_38_clk), .rst(icmp_38_rst),
		.data_in_bus({icmp_38_in2_data, icmp_38_in1_data}), .valid_in_bus({icmp_38_in2_valid, icmp_38_in1_valid}), .ready_in_bus({icmp_38_in2_ready, icmp_38_in1_ready}), 
		.data_out_bus({icmp_38_out1_data}), .valid_out_bus({icmp_38_out1_valid}), .ready_out_bus({icmp_38_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n0
		(.clk(phi_n0_clk), .rst(phi_n0_rst),
		.data_in_bus({phi_n0_in1_data}), .valid_in_bus({phi_n0_in1_valid}), .ready_in_bus({phi_n0_in1_ready}), 
		.data_out_bus({phi_n0_out1_data}), .valid_out_bus({phi_n0_out1_valid}), .ready_out_bus({phi_n0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n1
		(.clk(phi_n1_clk), .rst(phi_n1_rst),
		.data_in_bus({phi_n1_in1_data}), .valid_in_bus({phi_n1_in1_valid}), .ready_in_bus({phi_n1_in1_ready}), 
		.data_out_bus({phi_n1_out1_data}), .valid_out_bus({phi_n1_out1_valid}), .ready_out_bus({phi_n1_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_5
		(.clk(fork_5_clk), .rst(fork_5_rst),
		.data_in_bus({fork_5_in1_data}), .valid_in_bus({fork_5_in1_valid}), .ready_in_bus({fork_5_in1_ready}), 
		.data_out_bus({fork_5_out2_data, fork_5_out1_data}), .valid_out_bus({fork_5_out2_valid, fork_5_out1_valid}), .ready_out_bus({fork_5_out2_ready, fork_5_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_24
		(.clk(branch_24_clk), .rst(branch_24_rst),
		.data_in_bus({{31'b0, branch_24_in2_data}, branch_24_in1_data}), .valid_in_bus({branch_24_in2_valid, branch_24_in1_valid}), .ready_in_bus({branch_24_in2_ready, branch_24_in1_ready}), 
		.data_out_bus({branch_24_out2_data, branch_24_out1_data}), .valid_out_bus({branch_24_out2_valid, branch_24_out1_valid}), .ready_out_bus({branch_24_out2_ready, branch_24_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_25
		(.clk(branch_25_clk), .rst(branch_25_rst),
		.data_in_bus({{4'b0, branch_25_in2_data}, branch_25_in1_data}), .valid_in_bus({branch_25_in2_valid, branch_25_in1_valid}), .ready_in_bus({branch_25_in2_ready, branch_25_in1_ready}), 
		.data_out_bus({branch_25_out2_data, branch_25_out1_data}), .valid_out_bus({branch_25_out2_valid, branch_25_out1_valid}), .ready_out_bus({branch_25_out2_ready, branch_25_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_22
		(.clk(fork_22_clk), .rst(fork_22_rst),
		.data_in_bus({fork_22_in1_data}), .valid_in_bus({fork_22_in1_valid}), .ready_in_bus({fork_22_in1_ready}), 
		.data_out_bus({fork_22_out3_data, fork_22_out2_data, fork_22_out1_data}), .valid_out_bus({fork_22_out3_valid, fork_22_out2_valid, fork_22_out1_valid}), .ready_out_bus({fork_22_out3_ready, fork_22_out2_ready, fork_22_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_22
		(.clk(phiC_22_clk), .rst(phiC_22_rst),
		.data_in_bus({phiC_22_in1_data}), .valid_in_bus({phiC_22_in1_valid}), .ready_in_bus({phiC_22_in1_ready}), 
		.data_out_bus({phiC_22_out1_data}), .valid_out_bus({phiC_22_out1_valid}), .ready_out_bus({phiC_22_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_33
		(.clk(branchC_33_clk), .rst(branchC_33_rst),
		.data_in_bus({{branchC_33_in2_data}, branchC_33_in1_data}), .valid_in_bus({branchC_33_in2_valid, branchC_33_in1_valid}), .ready_in_bus({branchC_33_in2_ready, branchC_33_in1_ready}), 
		.data_out_bus({branchC_33_out2_data, branchC_33_out1_data}), .valid_out_bus({branchC_33_out2_valid, branchC_33_out1_valid}), .ready_out_bus({branchC_33_out2_ready, branchC_33_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_9
		(.clk(source_9_clk), .rst(source_9_rst),
		.data_out_bus({source_9_out1_data}), .valid_out_bus({source_9_out1_valid}), .ready_out_bus({source_9_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(5))source_node_source_10
		(.clk(source_10_clk), .rst(source_10_rst),
		.data_out_bus({source_10_out1_data}), .valid_out_bus({source_10_out1_valid}), .ready_out_bus({source_10_out1_ready}));

	ret_op #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) ret_op_ret_0
		(.clk(ret_0_clk), .rst(ret_0_rst),
		.data_in_bus({ret_0_in1_data}), .valid_in_bus({ret_0_in1_valid}), .ready_in_bus({ret_0_in1_ready}), 
		.data_out_bus({ret_0_out1_data}), .valid_out_bus({ret_0_out1_valid}), .ready_out_bus({ret_0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n15
		(.clk(phi_n15_clk), .rst(phi_n15_rst),
		.data_in_bus({phi_n15_in1_data}), .valid_in_bus({phi_n15_in1_valid}), .ready_in_bus({phi_n15_in1_ready}), 
		.data_out_bus({phi_n15_out1_data}), .valid_out_bus({phi_n15_out1_valid}), .ready_out_bus({phi_n15_out1_ready}));

	end_node #(.INPUTS(1), .OUTPUTS(1), .MEMORY_INPUTS(3), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) end_node_end_0
		(.clk(end_0_clk), .rst(end_0_rst),
		.data_in_bus({end_0_in4_data}), .valid_in_bus({end_0_in4_valid}), .ready_in_bus({end_0_in4_ready}), .e_valid_bus({end_0_in3_valid, end_0_in2_valid, end_0_in1_valid}), .e_ready_bus({end_0_in3_ready, end_0_in2_ready, end_0_in1_ready}), 
		.data_out_bus({end_0_out1_data}), .valid_out_bus({end_0_out1_valid}), .ready_out_bus({end_0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_23
		(.clk(phiC_23_clk), .rst(phiC_23_rst),
		.data_in_bus({phiC_23_in1_data}), .valid_in_bus({phiC_23_in1_valid}), .ready_in_bus({phiC_23_in1_ready}), 
		.data_out_bus({phiC_23_out1_data}), .valid_out_bus({phiC_23_out1_valid}), .ready_out_bus({phiC_23_out1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_0
		(.clk(sink_0_clk), .rst(sink_0_rst),
		.data_in_bus({sink_0_in1_data}), .valid_in_bus({sink_0_in1_valid}), .ready_in_bus({sink_0_in1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5), .COND_SIZE(1)) mux_node_phi_3
		(.clk(phi_3_clk), .rst(phi_3_rst),
		.data_in_bus({{4'b0, phi_3_in1_data}, phi_3_in3_data, phi_3_in2_data}), .valid_in_bus({phi_3_in1_valid, phi_3_in3_valid, phi_3_in2_valid}), .ready_in_bus({phi_3_in1_ready, phi_3_in3_ready, phi_3_in2_ready}), 
		.data_out_bus({phi_3_out1_data}), .valid_out_bus({phi_3_out1_valid}), .ready_out_bus({phi_3_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block3
		(.clk(brCst_block3_clk), .rst(brCst_block3_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block3_in1_valid}), .ready_in_bus({brCst_block3_in1_ready}), 
		.data_out_bus({brCst_block3_out1_data}), .valid_out_bus({brCst_block3_out1_valid}), .ready_out_bus({brCst_block3_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_2
		(.clk(cst_2_clk), .rst(cst_2_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_2_in1_valid}), .ready_in_bus({cst_2_in1_ready}), 
		.data_out_bus({cst_2_out1_data}), .valid_out_bus({cst_2_out1_valid}), .ready_out_bus({cst_2_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_3
		(.clk(cst_3_clk), .rst(cst_3_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_3_in1_valid}), .ready_in_bus({cst_3_in1_ready}), 
		.data_out_bus({cst_3_out1_data}), .valid_out_bus({cst_3_out1_valid}), .ready_out_bus({cst_3_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n2
		(.clk(phi_n2_clk), .rst(phi_n2_rst),
		.data_in_bus({phi_n2_in2_data, phi_n2_in1_data}), .valid_in_bus({phi_n2_in2_valid, phi_n2_in1_valid}), .ready_in_bus({phi_n2_in2_ready, phi_n2_in1_ready}), 
		.data_out_bus({phi_n2_out1_data}), .valid_out_bus({phi_n2_out1_valid}), .ready_out_bus({phi_n2_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_3
		(.clk(branch_3_clk), .rst(branch_3_rst),
		.data_in_bus({{branch_3_in2_data}, branch_3_in1_data}), .valid_in_bus({branch_3_in2_valid, branch_3_in1_valid}), .ready_in_bus({branch_3_in2_ready, branch_3_in1_ready}), 
		.data_out_bus({branch_3_out2_data, branch_3_out1_data}), .valid_out_bus({branch_3_out2_valid, branch_3_out1_valid}), .ready_out_bus({branch_3_out2_ready, branch_3_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_4
		(.clk(branch_4_clk), .rst(branch_4_rst),
		.data_in_bus({{branch_4_in2_data}, branch_4_in1_data}), .valid_in_bus({branch_4_in2_valid, branch_4_in1_valid}), .ready_in_bus({branch_4_in2_ready, branch_4_in1_ready}), 
		.data_out_bus({branch_4_out2_data, branch_4_out1_data}), .valid_out_bus({branch_4_out2_valid, branch_4_out1_valid}), .ready_out_bus({branch_4_out2_ready, branch_4_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_5
		(.clk(branch_5_clk), .rst(branch_5_rst),
		.data_in_bus({{4'b0, branch_5_in2_data}, branch_5_in1_data}), .valid_in_bus({branch_5_in2_valid, branch_5_in1_valid}), .ready_in_bus({branch_5_in2_ready, branch_5_in1_ready}), 
		.data_out_bus({branch_5_out2_data, branch_5_out1_data}), .valid_out_bus({branch_5_out2_valid, branch_5_out1_valid}), .ready_out_bus({branch_5_out2_ready, branch_5_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_6
		(.clk(branch_6_clk), .rst(branch_6_rst),
		.data_in_bus({{4'b0, branch_6_in2_data}, branch_6_in1_data}), .valid_in_bus({branch_6_in2_valid, branch_6_in1_valid}), .ready_in_bus({branch_6_in2_ready, branch_6_in1_ready}), 
		.data_out_bus({branch_6_out2_data, branch_6_out1_data}), .valid_out_bus({branch_6_out2_valid, branch_6_out1_valid}), .ready_out_bus({branch_6_out2_ready, branch_6_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_17
		(.clk(fork_17_clk), .rst(fork_17_rst),
		.data_in_bus({fork_17_in1_data}), .valid_in_bus({fork_17_in1_valid}), .ready_in_bus({fork_17_in1_ready}), 
		.data_out_bus({fork_17_out5_data, fork_17_out4_data, fork_17_out3_data, fork_17_out2_data, fork_17_out1_data}), .valid_out_bus({fork_17_out5_valid, fork_17_out4_valid, fork_17_out3_valid, fork_17_out2_valid, fork_17_out1_valid}), .ready_out_bus({fork_17_out5_ready, fork_17_out4_ready, fork_17_out3_ready, fork_17_out2_ready, fork_17_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_17
		(.clk(phiC_17_clk), .rst(phiC_17_rst),
		.data_in_bus({phiC_17_in2_data, phiC_17_in1_data}), .valid_in_bus({phiC_17_in2_valid, phiC_17_in1_valid}), .ready_in_bus({phiC_17_in2_ready, phiC_17_in1_ready}), 
		.data_out_bus({phiC_17_out2_data, phiC_17_out1_data}), .valid_out_bus({phiC_17_out2_valid, phiC_17_out1_valid}), .ready_out_bus({phiC_17_out2_ready, phiC_17_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_27
		(.clk(forkC_27_clk), .rst(forkC_27_rst),
		.data_in_bus({forkC_27_in1_data}), .valid_in_bus({forkC_27_in1_valid}), .ready_in_bus({forkC_27_in1_ready}), 
		.data_out_bus({forkC_27_out4_data, forkC_27_out3_data, forkC_27_out2_data, forkC_27_out1_data}), .valid_out_bus({forkC_27_out4_valid, forkC_27_out3_valid, forkC_27_out2_valid, forkC_27_out1_valid}), .ready_out_bus({forkC_27_out4_ready, forkC_27_out3_ready, forkC_27_out2_ready, forkC_27_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_28
		(.clk(branchC_28_clk), .rst(branchC_28_rst),
		.data_in_bus({{branchC_28_in2_data}, branchC_28_in1_data}), .valid_in_bus({branchC_28_in2_valid, branchC_28_in1_valid}), .ready_in_bus({branchC_28_in2_ready, branchC_28_in1_ready}), 
		.data_out_bus({branchC_28_out2_data, branchC_28_out1_data}), .valid_out_bus({branchC_28_out2_valid, branchC_28_out1_valid}), .ready_out_bus({branchC_28_out2_ready, branchC_28_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) const_node_cst_11
		(.clk(cst_11_clk), .rst(cst_11_rst),
		.data_in_bus({5'd30}), .valid_in_bus({cst_11_in1_valid}), .ready_in_bus({cst_11_in1_ready}), 
		.data_out_bus({cst_11_out1_data}), .valid_out_bus({cst_11_out1_valid}), .ready_out_bus({cst_11_out1_ready}));

	mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(10)) mul_op_mul_30
		(.clk(mul_30_clk), .rst(mul_30_rst),
		.data_in_bus({mul_30_in2_data, mul_30_in1_data}), .valid_in_bus({mul_30_in2_valid, mul_30_in1_valid}), .ready_in_bus({mul_30_in2_ready, mul_30_in1_ready}), 
		.data_out_bus({mul_30_out1_data}), .valid_out_bus({mul_30_out1_valid}), .ready_out_bus({mul_30_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(11), .DATA_OUT_SIZE(11)) add_op_add_31
		(.clk(add_31_clk), .rst(add_31_rst),
		.data_in_bus({add_31_in2_data, add_31_in1_data}), .valid_in_bus({add_31_in2_valid, add_31_in1_valid}), .ready_in_bus({add_31_in2_ready, add_31_in1_ready}), 
		.data_out_bus({add_31_out1_data}), .valid_out_bus({add_31_out1_valid}), .ready_out_bus({add_31_out1_ready}));

	mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(11), .DATA_SIZE(32)) mc_store_op_store_0
		(.clk(store_0_clk), .rst(store_0_rst),
		.data_in_bus({store_0_in1_data}), .address_in_bus({store_0_in2_data}), .valid_in_bus({store_0_in2_valid, store_0_in1_valid}), .ready_in_bus({store_0_in2_ready, store_0_in1_ready}), 
		.data_out_bus({store_0_out1_data}), .address_out_bus({store_0_out2_data}), .valid_out_bus({store_0_out2_valid, store_0_out1_valid}), .ready_out_bus({store_0_out2_ready, store_0_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_12
		(.clk(cst_12_clk), .rst(cst_12_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_12_in1_valid}), .ready_in_bus({cst_12_in1_ready}), 
		.data_out_bus({cst_12_out1_data}), .valid_out_bus({cst_12_out1_valid}), .ready_out_bus({cst_12_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) add_op_add_34
		(.clk(add_34_clk), .rst(add_34_rst),
		.data_in_bus({add_34_in2_data, add_34_in1_data}), .valid_in_bus({add_34_in2_valid, add_34_in1_valid}), .ready_in_bus({add_34_in2_ready, add_34_in1_ready}), 
		.data_out_bus({add_34_out1_data}), .valid_out_bus({add_34_out1_valid}), .ready_out_bus({add_34_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) const_node_cst_13
		(.clk(cst_13_clk), .rst(cst_13_rst),
		.data_in_bus({5'd28}), .valid_in_bus({cst_13_in1_valid}), .ready_in_bus({cst_13_in1_ready}), 
		.data_out_bus({cst_13_out1_data}), .valid_out_bus({cst_13_out1_valid}), .ready_out_bus({cst_13_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_35
		(.clk(icmp_35_clk), .rst(icmp_35_rst),
		.data_in_bus({icmp_35_in2_data, icmp_35_in1_data}), .valid_in_bus({icmp_35_in2_valid, icmp_35_in1_valid}), .ready_in_bus({icmp_35_in2_ready, icmp_35_in1_ready}), 
		.data_out_bus({icmp_35_out1_data}), .valid_out_bus({icmp_35_out1_valid}), .ready_out_bus({icmp_35_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n3
		(.clk(phi_n3_clk), .rst(phi_n3_rst),
		.data_in_bus({phi_n3_in1_data}), .valid_in_bus({phi_n3_in1_valid}), .ready_in_bus({phi_n3_in1_ready}), 
		.data_out_bus({phi_n3_out1_data}), .valid_out_bus({phi_n3_out1_valid}), .ready_out_bus({phi_n3_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n4
		(.clk(phi_n4_clk), .rst(phi_n4_rst),
		.data_in_bus({phi_n4_in1_data}), .valid_in_bus({phi_n4_in1_valid}), .ready_in_bus({phi_n4_in1_ready}), 
		.data_out_bus({phi_n4_out1_data}), .valid_out_bus({phi_n4_out1_valid}), .ready_out_bus({phi_n4_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n5
		(.clk(phi_n5_clk), .rst(phi_n5_rst),
		.data_in_bus({phi_n5_in1_data}), .valid_in_bus({phi_n5_in1_valid}), .ready_in_bus({phi_n5_in1_ready}), 
		.data_out_bus({phi_n5_out1_data}), .valid_out_bus({phi_n5_out1_valid}), .ready_out_bus({phi_n5_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_4
		(.clk(fork_4_clk), .rst(fork_4_rst),
		.data_in_bus({fork_4_in1_data}), .valid_in_bus({fork_4_in1_valid}), .ready_in_bus({fork_4_in1_ready}), 
		.data_out_bus({fork_4_out2_data, fork_4_out1_data}), .valid_out_bus({fork_4_out2_valid, fork_4_out1_valid}), .ready_out_bus({fork_4_out2_ready, fork_4_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_6
		(.clk(fork_6_clk), .rst(fork_6_rst),
		.data_in_bus({fork_6_in1_data}), .valid_in_bus({fork_6_in1_valid}), .ready_in_bus({fork_6_in1_ready}), 
		.data_out_bus({fork_6_out2_data, fork_6_out1_data}), .valid_out_bus({fork_6_out2_valid, fork_6_out1_valid}), .ready_out_bus({fork_6_out2_ready, fork_6_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_7
		(.clk(fork_7_clk), .rst(fork_7_rst),
		.data_in_bus({fork_7_in1_data}), .valid_in_bus({fork_7_in1_valid}), .ready_in_bus({fork_7_in1_ready}), 
		.data_out_bus({fork_7_out2_data, fork_7_out1_data}), .valid_out_bus({fork_7_out2_valid, fork_7_out1_valid}), .ready_out_bus({fork_7_out2_ready, fork_7_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_8
		(.clk(fork_8_clk), .rst(fork_8_rst),
		.data_in_bus({fork_8_in1_data}), .valid_in_bus({fork_8_in1_valid}), .ready_in_bus({fork_8_in1_ready}), 
		.data_out_bus({fork_8_out2_data, fork_8_out1_data}), .valid_out_bus({fork_8_out2_valid, fork_8_out1_valid}), .ready_out_bus({fork_8_out2_ready, fork_8_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_21
		(.clk(branch_21_clk), .rst(branch_21_rst),
		.data_in_bus({{4'b0, branch_21_in2_data}, branch_21_in1_data}), .valid_in_bus({branch_21_in2_valid, branch_21_in1_valid}), .ready_in_bus({branch_21_in2_ready, branch_21_in1_ready}), 
		.data_out_bus({branch_21_out2_data, branch_21_out1_data}), .valid_out_bus({branch_21_out2_valid, branch_21_out1_valid}), .ready_out_bus({branch_21_out2_ready, branch_21_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_22
		(.clk(branch_22_clk), .rst(branch_22_rst),
		.data_in_bus({{4'b0, branch_22_in2_data}, branch_22_in1_data}), .valid_in_bus({branch_22_in2_valid, branch_22_in1_valid}), .ready_in_bus({branch_22_in2_ready, branch_22_in1_ready}), 
		.data_out_bus({branch_22_out2_data, branch_22_out1_data}), .valid_out_bus({branch_22_out2_valid, branch_22_out1_valid}), .ready_out_bus({branch_22_out2_ready, branch_22_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_23
		(.clk(branch_23_clk), .rst(branch_23_rst),
		.data_in_bus({{31'b0, branch_23_in2_data}, branch_23_in1_data}), .valid_in_bus({branch_23_in2_valid, branch_23_in1_valid}), .ready_in_bus({branch_23_in2_ready, branch_23_in1_ready}), 
		.data_out_bus({branch_23_out2_data, branch_23_out1_data}), .valid_out_bus({branch_23_out2_valid, branch_23_out1_valid}), .ready_out_bus({branch_23_out2_ready, branch_23_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_21
		(.clk(fork_21_clk), .rst(fork_21_rst),
		.data_in_bus({fork_21_in1_data}), .valid_in_bus({fork_21_in1_valid}), .ready_in_bus({fork_21_in1_ready}), 
		.data_out_bus({fork_21_out4_data, fork_21_out3_data, fork_21_out2_data, fork_21_out1_data}), .valid_out_bus({fork_21_out4_valid, fork_21_out3_valid, fork_21_out2_valid, fork_21_out1_valid}), .ready_out_bus({fork_21_out4_ready, fork_21_out3_ready, fork_21_out2_ready, fork_21_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_16
		(.clk(cst_16_clk), .rst(cst_16_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_16_in1_valid}), .ready_in_bus({cst_16_in1_ready}), 
		.data_out_bus({cst_16_out1_data}), .valid_out_bus({cst_16_out1_valid}), .ready_out_bus({cst_16_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_21
		(.clk(phiC_21_clk), .rst(phiC_21_rst),
		.data_in_bus({phiC_21_in1_data}), .valid_in_bus({phiC_21_in1_valid}), .ready_in_bus({phiC_21_in1_ready}), 
		.data_out_bus({phiC_21_out1_data}), .valid_out_bus({phiC_21_out1_valid}), .ready_out_bus({phiC_21_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_31
		(.clk(forkC_31_clk), .rst(forkC_31_rst),
		.data_in_bus({forkC_31_in1_data}), .valid_in_bus({forkC_31_in1_valid}), .ready_in_bus({forkC_31_in1_ready}), 
		.data_out_bus({forkC_31_out2_data, forkC_31_out1_data}), .valid_out_bus({forkC_31_out2_valid, forkC_31_out1_valid}), .ready_out_bus({forkC_31_out2_ready, forkC_31_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_32
		(.clk(branchC_32_clk), .rst(branchC_32_rst),
		.data_in_bus({{branchC_32_in2_data}, branchC_32_in1_data}), .valid_in_bus({branchC_32_in2_valid, branchC_32_in1_valid}), .ready_in_bus({branchC_32_in2_ready, branchC_32_in1_ready}), 
		.data_out_bus({branchC_32_out2_data, branchC_32_out1_data}), .valid_out_bus({branchC_32_out2_valid, branchC_32_out1_valid}), .ready_out_bus({branchC_32_out2_ready, branchC_32_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(5))source_node_source_6
		(.clk(source_6_clk), .rst(source_6_rst),
		.data_out_bus({source_6_out1_data}), .valid_out_bus({source_6_out1_valid}), .ready_out_bus({source_6_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_7
		(.clk(source_7_clk), .rst(source_7_rst),
		.data_out_bus({source_7_out1_data}), .valid_out_bus({source_7_out1_valid}), .ready_out_bus({source_7_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(5))source_node_source_8
		(.clk(source_8_clk), .rst(source_8_rst),
		.data_out_bus({source_8_out1_data}), .valid_out_bus({source_8_out1_valid}), .ready_out_bus({source_8_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5), .COND_SIZE(1)) mux_node_phi_1
		(.clk(phi_1_clk), .rst(phi_1_rst),
		.data_in_bus({{4'b0, phi_1_in1_data}, phi_1_in3_data, phi_1_in2_data}), .valid_in_bus({phi_1_in1_valid, phi_1_in3_valid, phi_1_in2_valid}), .ready_in_bus({phi_1_in1_ready, phi_1_in3_ready, phi_1_in2_ready}), 
		.data_out_bus({phi_1_out1_data}), .valid_out_bus({phi_1_out1_valid}), .ready_out_bus({phi_1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block2
		(.clk(brCst_block2_clk), .rst(brCst_block2_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block2_in1_valid}), .ready_in_bus({brCst_block2_in1_ready}), 
		.data_out_bus({brCst_block2_out1_data}), .valid_out_bus({brCst_block2_out1_valid}), .ready_out_bus({brCst_block2_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_1
		(.clk(cst_1_clk), .rst(cst_1_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_1_in1_valid}), .ready_in_bus({cst_1_in1_ready}), 
		.data_out_bus({cst_1_out1_data}), .valid_out_bus({cst_1_out1_valid}), .ready_out_bus({cst_1_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_1
		(.clk(branch_1_clk), .rst(branch_1_rst),
		.data_in_bus({{branch_1_in2_data}, branch_1_in1_data}), .valid_in_bus({branch_1_in2_valid, branch_1_in1_valid}), .ready_in_bus({branch_1_in2_ready, branch_1_in1_ready}), 
		.data_out_bus({branch_1_out2_data, branch_1_out1_data}), .valid_out_bus({branch_1_out2_valid, branch_1_out1_valid}), .ready_out_bus({branch_1_out2_ready, branch_1_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_2
		(.clk(branch_2_clk), .rst(branch_2_rst),
		.data_in_bus({{4'b0, branch_2_in2_data}, branch_2_in1_data}), .valid_in_bus({branch_2_in2_valid, branch_2_in1_valid}), .ready_in_bus({branch_2_in2_ready, branch_2_in1_ready}), 
		.data_out_bus({branch_2_out2_data, branch_2_out1_data}), .valid_out_bus({branch_2_out2_valid, branch_2_out1_valid}), .ready_out_bus({branch_2_out2_ready, branch_2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_16
		(.clk(fork_16_clk), .rst(fork_16_rst),
		.data_in_bus({fork_16_in1_data}), .valid_in_bus({fork_16_in1_valid}), .ready_in_bus({fork_16_in1_ready}), 
		.data_out_bus({fork_16_out3_data, fork_16_out2_data, fork_16_out1_data}), .valid_out_bus({fork_16_out3_valid, fork_16_out2_valid, fork_16_out1_valid}), .ready_out_bus({fork_16_out3_ready, fork_16_out2_ready, fork_16_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_16
		(.clk(phiC_16_clk), .rst(phiC_16_rst),
		.data_in_bus({phiC_16_in2_data, phiC_16_in1_data}), .valid_in_bus({phiC_16_in2_valid, phiC_16_in1_valid}), .ready_in_bus({phiC_16_in2_ready, phiC_16_in1_ready}), 
		.data_out_bus({phiC_16_out2_data, phiC_16_out1_data}), .valid_out_bus({phiC_16_out2_valid, phiC_16_out1_valid}), .ready_out_bus({phiC_16_out2_ready, phiC_16_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_26
		(.clk(forkC_26_clk), .rst(forkC_26_rst),
		.data_in_bus({forkC_26_in1_data}), .valid_in_bus({forkC_26_in1_valid}), .ready_in_bus({forkC_26_in1_ready}), 
		.data_out_bus({forkC_26_out3_data, forkC_26_out2_data, forkC_26_out1_data}), .valid_out_bus({forkC_26_out3_valid, forkC_26_out2_valid, forkC_26_out1_valid}), .ready_out_bus({forkC_26_out3_ready, forkC_26_out2_ready, forkC_26_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_27
		(.clk(branchC_27_clk), .rst(branchC_27_rst),
		.data_in_bus({{branchC_27_in2_data}, branchC_27_in1_data}), .valid_in_bus({branchC_27_in2_valid, branchC_27_in1_valid}), .ready_in_bus({branchC_27_in2_ready, branchC_27_in1_ready}), 
		.data_out_bus({branchC_27_out2_data, branchC_27_out1_data}), .valid_out_bus({branchC_27_out2_valid, branchC_27_out1_valid}), .ready_out_bus({branchC_27_out2_ready, branchC_27_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3), .COND_SIZE(1)) mux_node_phi_8
		(.clk(phi_8_clk), .rst(phi_8_rst),
		.data_in_bus({{2'b0, phi_8_in1_data}, phi_8_in3_data, phi_8_in2_data}), .valid_in_bus({phi_8_in1_valid, phi_8_in3_valid, phi_8_in2_valid}), .ready_in_bus({phi_8_in1_ready, phi_8_in3_ready, phi_8_in2_ready}), 
		.data_out_bus({phi_8_out1_data}), .valid_out_bus({phi_8_out1_valid}), .ready_out_bus({phi_8_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_9
		(.clk(phi_9_clk), .rst(phi_9_rst),
		.data_in_bus({{31'b0, phi_9_in1_data}, phi_9_in3_data, phi_9_in2_data}), .valid_in_bus({phi_9_in1_valid, phi_9_in3_valid, phi_9_in2_valid}), .ready_in_bus({phi_9_in1_ready, phi_9_in3_ready, phi_9_in2_ready}), 
		.data_out_bus({phi_9_out1_data}), .valid_out_bus({phi_9_out1_valid}), .ready_out_bus({phi_9_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_5
		(.clk(cst_5_clk), .rst(cst_5_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_5_in1_valid}), .ready_in_bus({cst_5_in1_ready}), 
		.data_out_bus({cst_5_out1_data}), .valid_out_bus({cst_5_out1_valid}), .ready_out_bus({cst_5_out1_ready}));

	mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(5)) mul_op_mul_10
		(.clk(mul_10_clk), .rst(mul_10_rst),
		.data_in_bus({mul_10_in2_data, mul_10_in1_data}), .valid_in_bus({mul_10_in2_valid, mul_10_in1_valid}), .ready_in_bus({mul_10_in2_ready, mul_10_in1_ready}), 
		.data_out_bus({mul_10_out1_data}), .valid_out_bus({mul_10_out1_valid}), .ready_out_bus({mul_10_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_11
		(.clk(add_11_clk), .rst(add_11_rst),
		.data_in_bus({add_11_in2_data, add_11_in1_data}), .valid_in_bus({add_11_in2_valid, add_11_in1_valid}), .ready_in_bus({add_11_in2_ready, add_11_in1_ready}), 
		.data_out_bus({add_11_out1_data}), .valid_out_bus({add_11_out1_valid}), .ready_out_bus({add_11_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(6), .DATA_SIZE(32)) mc_load_op_load_14
		(.clk(load_14_clk), .rst(load_14_rst),
		.data_in_bus({load_14_in1_data}), .address_in_bus({load_14_in2_data}), .valid_in_bus({load_14_in2_valid, load_14_in1_valid}), .ready_in_bus({load_14_in2_ready, load_14_in1_ready}), 
		.data_out_bus({load_14_out1_data}), .address_out_bus({load_14_out2_data}), .valid_out_bus({load_14_out2_valid, load_14_out1_valid}), .ready_out_bus({load_14_out2_ready, load_14_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_15
		(.clk(add_15_clk), .rst(add_15_rst),
		.data_in_bus({add_15_in2_data, add_15_in1_data}), .valid_in_bus({add_15_in2_valid, add_15_in1_valid}), .ready_in_bus({add_15_in2_ready, add_15_in1_ready}), 
		.data_out_bus({add_15_out1_data}), .valid_out_bus({add_15_out1_valid}), .ready_out_bus({add_15_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) const_node_cst_6
		(.clk(cst_6_clk), .rst(cst_6_rst),
		.data_in_bus({5'd30}), .valid_in_bus({cst_6_in1_valid}), .ready_in_bus({cst_6_in1_ready}), 
		.data_out_bus({cst_6_out1_data}), .valid_out_bus({cst_6_out1_valid}), .ready_out_bus({cst_6_out1_ready}));

	mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(11)) mul_op_mul_16
		(.clk(mul_16_clk), .rst(mul_16_rst),
		.data_in_bus({mul_16_in2_data, mul_16_in1_data}), .valid_in_bus({mul_16_in2_valid, mul_16_in1_valid}), .ready_in_bus({mul_16_in2_ready, mul_16_in1_ready}), 
		.data_out_bus({mul_16_out1_data}), .valid_out_bus({mul_16_out1_valid}), .ready_out_bus({mul_16_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(12), .DATA_OUT_SIZE(12)) add_op_add_17
		(.clk(add_17_clk), .rst(add_17_rst),
		.data_in_bus({add_17_in2_data, add_17_in1_data}), .valid_in_bus({add_17_in2_valid, add_17_in1_valid}), .ready_in_bus({add_17_in2_ready, add_17_in1_ready}), 
		.data_out_bus({add_17_out1_data}), .valid_out_bus({add_17_out1_valid}), .ready_out_bus({add_17_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(13), .DATA_OUT_SIZE(13)) add_op_add_18
		(.clk(add_18_clk), .rst(add_18_rst),
		.data_in_bus({add_18_in2_data, add_18_in1_data}), .valid_in_bus({add_18_in2_valid, add_18_in1_valid}), .ready_in_bus({add_18_in2_ready, add_18_in1_ready}), 
		.data_out_bus({add_18_out1_data}), .valid_out_bus({add_18_out1_valid}), .ready_out_bus({add_18_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(13), .DATA_SIZE(32)) mc_load_op_load_21
		(.clk(load_21_clk), .rst(load_21_rst),
		.data_in_bus({load_21_in1_data}), .address_in_bus({load_21_in2_data}), .valid_in_bus({load_21_in2_valid, load_21_in1_valid}), .ready_in_bus({load_21_in2_ready, load_21_in1_ready}), 
		.data_out_bus({load_21_out1_data}), .address_out_bus({load_21_out2_data}), .valid_out_bus({load_21_out2_valid, load_21_out1_valid}), .ready_out_bus({load_21_out2_ready, load_21_out1_ready}));

	mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(16), .DATA_OUT_SIZE(32)) mul_op_mul_22
		(.clk(mul_22_clk), .rst(mul_22_rst),
		.data_in_bus({mul_22_in2_data, mul_22_in1_data}), .valid_in_bus({mul_22_in2_valid, mul_22_in1_valid}), .ready_in_bus({mul_22_in2_ready, mul_22_in1_ready}), 
		.data_out_bus({mul_22_out1_data}), .valid_out_bus({mul_22_out1_valid}), .ready_out_bus({mul_22_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_23
		(.clk(add_23_clk), .rst(add_23_rst),
		.data_in_bus({add_23_in2_data, add_23_in1_data}), .valid_in_bus({add_23_in2_valid, add_23_in1_valid}), .ready_in_bus({add_23_in2_ready, add_23_in1_ready}), 
		.data_out_bus({add_23_out1_data}), .valid_out_bus({add_23_out1_valid}), .ready_out_bus({add_23_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_7
		(.clk(cst_7_clk), .rst(cst_7_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_7_in1_valid}), .ready_in_bus({cst_7_in1_ready}), 
		.data_out_bus({cst_7_out1_data}), .valid_out_bus({cst_7_out1_valid}), .ready_out_bus({cst_7_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) add_op_add_24
		(.clk(add_24_clk), .rst(add_24_rst),
		.data_in_bus({add_24_in2_data, add_24_in1_data}), .valid_in_bus({add_24_in2_valid, add_24_in1_valid}), .ready_in_bus({add_24_in2_ready, add_24_in1_ready}), 
		.data_out_bus({add_24_out1_data}), .valid_out_bus({add_24_out1_valid}), .ready_out_bus({add_24_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_8
		(.clk(cst_8_clk), .rst(cst_8_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_8_in1_valid}), .ready_in_bus({cst_8_in1_ready}), 
		.data_out_bus({cst_8_out1_data}), .valid_out_bus({cst_8_out1_valid}), .ready_out_bus({cst_8_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_25
		(.clk(icmp_25_clk), .rst(icmp_25_rst),
		.data_in_bus({icmp_25_in2_data, icmp_25_in1_data}), .valid_in_bus({icmp_25_in2_valid, icmp_25_in1_valid}), .ready_in_bus({icmp_25_in2_ready, icmp_25_in1_ready}), 
		.data_out_bus({icmp_25_out1_data}), .valid_out_bus({icmp_25_out1_valid}), .ready_out_bus({icmp_25_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) merge_node_phi_n12
		(.clk(phi_n12_clk), .rst(phi_n12_rst),
		.data_in_bus({phi_n12_in2_data, phi_n12_in1_data}), .valid_in_bus({phi_n12_in2_valid, phi_n12_in1_valid}), .ready_in_bus({phi_n12_in2_ready, phi_n12_in1_ready}), 
		.data_out_bus({phi_n12_out1_data}), .valid_out_bus({phi_n12_out1_valid}), .ready_out_bus({phi_n12_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n13
		(.clk(phi_n13_clk), .rst(phi_n13_rst),
		.data_in_bus({phi_n13_in2_data, phi_n13_in1_data}), .valid_in_bus({phi_n13_in2_valid, phi_n13_in1_valid}), .ready_in_bus({phi_n13_in2_ready, phi_n13_in1_ready}), 
		.data_out_bus({phi_n13_out1_data}), .valid_out_bus({phi_n13_out1_valid}), .ready_out_bus({phi_n13_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) merge_node_phi_n14
		(.clk(phi_n14_clk), .rst(phi_n14_rst),
		.data_in_bus({phi_n14_in2_data, phi_n14_in1_data}), .valid_in_bus({phi_n14_in2_valid, phi_n14_in1_valid}), .ready_in_bus({phi_n14_in2_ready, phi_n14_in1_ready}), 
		.data_out_bus({phi_n14_out1_data}), .valid_out_bus({phi_n14_out1_valid}), .ready_out_bus({phi_n14_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) fork_node_fork_0
		(.clk(fork_0_clk), .rst(fork_0_rst),
		.data_in_bus({fork_0_in1_data}), .valid_in_bus({fork_0_in1_valid}), .ready_in_bus({fork_0_in1_ready}), 
		.data_out_bus({fork_0_out3_data, fork_0_out2_data, fork_0_out1_data}), .valid_out_bus({fork_0_out3_valid, fork_0_out2_valid, fork_0_out1_valid}), .ready_out_bus({fork_0_out3_ready, fork_0_out2_ready, fork_0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) fork_node_fork_2
		(.clk(fork_2_clk), .rst(fork_2_rst),
		.data_in_bus({fork_2_in1_data}), .valid_in_bus({fork_2_in1_valid}), .ready_in_bus({fork_2_in1_ready}), 
		.data_out_bus({fork_2_out2_data, fork_2_out1_data}), .valid_out_bus({fork_2_out2_valid, fork_2_out1_valid}), .ready_out_bus({fork_2_out2_ready, fork_2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) fork_node_fork_12
		(.clk(fork_12_clk), .rst(fork_12_rst),
		.data_in_bus({fork_12_in1_data}), .valid_in_bus({fork_12_in1_valid}), .ready_in_bus({fork_12_in1_ready}), 
		.data_out_bus({fork_12_out3_data, fork_12_out2_data, fork_12_out1_data}), .valid_out_bus({fork_12_out3_valid, fork_12_out2_valid, fork_12_out1_valid}), .ready_out_bus({fork_12_out3_ready, fork_12_out2_ready, fork_12_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_13
		(.clk(fork_13_clk), .rst(fork_13_rst),
		.data_in_bus({fork_13_in1_data}), .valid_in_bus({fork_13_in1_valid}), .ready_in_bus({fork_13_in1_ready}), 
		.data_out_bus({fork_13_out2_data, fork_13_out1_data}), .valid_out_bus({fork_13_out2_valid, fork_13_out1_valid}), .ready_out_bus({fork_13_out2_ready, fork_13_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) fork_node_fork_14
		(.clk(fork_14_clk), .rst(fork_14_rst),
		.data_in_bus({fork_14_in1_data}), .valid_in_bus({fork_14_in1_valid}), .ready_in_bus({fork_14_in1_ready}), 
		.data_out_bus({fork_14_out2_data, fork_14_out1_data}), .valid_out_bus({fork_14_out2_valid, fork_14_out1_valid}), .ready_out_bus({fork_14_out2_ready, fork_14_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_12
		(.clk(branch_12_clk), .rst(branch_12_rst),
		.data_in_bus({{31'b0, branch_12_in2_data}, branch_12_in1_data}), .valid_in_bus({branch_12_in2_valid, branch_12_in1_valid}), .ready_in_bus({branch_12_in2_ready, branch_12_in1_ready}), 
		.data_out_bus({branch_12_out2_data, branch_12_out1_data}), .valid_out_bus({branch_12_out2_valid, branch_12_out1_valid}), .ready_out_bus({branch_12_out2_ready, branch_12_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) branch_node_branch_13
		(.clk(branch_13_clk), .rst(branch_13_rst),
		.data_in_bus({{2'b0, branch_13_in2_data}, branch_13_in1_data}), .valid_in_bus({branch_13_in2_valid, branch_13_in1_valid}), .ready_in_bus({branch_13_in2_ready, branch_13_in1_ready}), 
		.data_out_bus({branch_13_out2_data, branch_13_out1_data}), .valid_out_bus({branch_13_out2_valid, branch_13_out1_valid}), .ready_out_bus({branch_13_out2_ready, branch_13_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) branch_node_branch_14
		(.clk(branch_14_clk), .rst(branch_14_rst),
		.data_in_bus({{2'b0, branch_14_in2_data}, branch_14_in1_data}), .valid_in_bus({branch_14_in2_valid, branch_14_in1_valid}), .ready_in_bus({branch_14_in2_ready, branch_14_in1_ready}), 
		.data_out_bus({branch_14_out2_data, branch_14_out1_data}), .valid_out_bus({branch_14_out2_valid, branch_14_out1_valid}), .ready_out_bus({branch_14_out2_ready, branch_14_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_15
		(.clk(branch_15_clk), .rst(branch_15_rst),
		.data_in_bus({{4'b0, branch_15_in2_data}, branch_15_in1_data}), .valid_in_bus({branch_15_in2_valid, branch_15_in1_valid}), .ready_in_bus({branch_15_in2_ready, branch_15_in1_ready}), 
		.data_out_bus({branch_15_out2_data, branch_15_out1_data}), .valid_out_bus({branch_15_out2_valid, branch_15_out1_valid}), .ready_out_bus({branch_15_out2_ready, branch_15_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(5), .DATA_OUT_SIZE(5)) branch_node_branch_16
		(.clk(branch_16_clk), .rst(branch_16_rst),
		.data_in_bus({{4'b0, branch_16_in2_data}, branch_16_in1_data}), .valid_in_bus({branch_16_in2_valid, branch_16_in1_valid}), .ready_in_bus({branch_16_in2_ready, branch_16_in1_ready}), 
		.data_out_bus({branch_16_out2_data, branch_16_out1_data}), .valid_out_bus({branch_16_out2_valid, branch_16_out1_valid}), .ready_out_bus({branch_16_out2_ready, branch_16_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(6), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_19
		(.clk(fork_19_clk), .rst(fork_19_rst),
		.data_in_bus({fork_19_in1_data}), .valid_in_bus({fork_19_in1_valid}), .ready_in_bus({fork_19_in1_ready}), 
		.data_out_bus({fork_19_out6_data, fork_19_out5_data, fork_19_out4_data, fork_19_out3_data, fork_19_out2_data, fork_19_out1_data}), .valid_out_bus({fork_19_out6_valid, fork_19_out5_valid, fork_19_out4_valid, fork_19_out3_valid, fork_19_out2_valid, fork_19_out1_valid}), .ready_out_bus({fork_19_out6_ready, fork_19_out5_ready, fork_19_out4_ready, fork_19_out3_ready, fork_19_out2_ready, fork_19_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_19
		(.clk(phiC_19_clk), .rst(phiC_19_rst),
		.data_in_bus({phiC_19_in2_data, phiC_19_in1_data}), .valid_in_bus({phiC_19_in2_valid, phiC_19_in1_valid}), .ready_in_bus({phiC_19_in2_ready, phiC_19_in1_ready}), 
		.data_out_bus({phiC_19_out2_data, phiC_19_out1_data}), .valid_out_bus({phiC_19_out2_valid, phiC_19_out1_valid}), .ready_out_bus({phiC_19_out2_ready, phiC_19_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_30
		(.clk(branchC_30_clk), .rst(branchC_30_rst),
		.data_in_bus({{branchC_30_in2_data}, branchC_30_in1_data}), .valid_in_bus({branchC_30_in2_valid, branchC_30_in1_valid}), .ready_in_bus({branchC_30_in2_ready, branchC_30_in1_ready}), 
		.data_out_bus({branchC_30_out2_data, branchC_30_out1_data}), .valid_out_bus({branchC_30_out2_valid, branchC_30_out1_valid}), .ready_out_bus({branchC_30_out2_ready, branchC_30_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_0
		(.clk(source_0_clk), .rst(source_0_rst),
		.data_out_bus({source_0_out1_data}), .valid_out_bus({source_0_out1_valid}), .ready_out_bus({source_0_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(5))source_node_source_1
		(.clk(source_1_clk), .rst(source_1_rst),
		.data_out_bus({source_1_out1_data}), .valid_out_bus({source_1_out1_valid}), .ready_out_bus({source_1_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_2
		(.clk(source_2_clk), .rst(source_2_rst),
		.data_out_bus({source_2_out1_data}), .valid_out_bus({source_2_out1_valid}), .ready_out_bus({source_2_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_3
		(.clk(source_3_clk), .rst(source_3_rst),
		.data_out_bus({source_3_out1_data}), .valid_out_bus({source_3_out1_valid}), .ready_out_bus({source_3_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_37
		(.clk(fork_37_clk), .rst(fork_37_rst),
		.data_in_bus({fork_37_in1_data}), .valid_in_bus({fork_37_in1_valid}), .ready_in_bus({fork_37_in1_ready}), 
		.data_out_bus({fork_37_out2_data, fork_37_out1_data}), .valid_out_bus({fork_37_out2_valid, fork_37_out1_valid}), .ready_out_bus({fork_37_out2_ready, fork_37_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block1
		(.clk(brCst_block1_clk), .rst(brCst_block1_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block1_in1_valid}), .ready_in_bus({brCst_block1_in1_ready}), 
		.data_out_bus({brCst_block1_out1_data}), .valid_out_bus({brCst_block1_out1_valid}), .ready_out_bus({brCst_block1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_0
		(.clk(cst_0_clk), .rst(cst_0_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_0_in1_valid}), .ready_in_bus({cst_0_in1_ready}), 
		.data_out_bus({cst_0_out1_data}), .valid_out_bus({cst_0_out1_valid}), .ready_out_bus({cst_0_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_0
		(.clk(branch_0_clk), .rst(branch_0_rst),
		.data_in_bus({{branch_0_in2_data}, branch_0_in1_data}), .valid_in_bus({branch_0_in2_valid, branch_0_in1_valid}), .ready_in_bus({branch_0_in2_ready, branch_0_in1_ready}), 
		.data_out_bus({branch_0_out2_data, branch_0_out1_data}), .valid_out_bus({branch_0_out2_valid, branch_0_out1_valid}), .ready_out_bus({branch_0_out2_ready, branch_0_out1_ready}));

	start_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) start_node_start_0
		(.clk(start_0_clk), .rst(start_0_rst),
		.data_in_bus({start_0_in1_data}), .valid_in_bus({start_0_in1_valid}), .ready_in_bus({start_0_in1_ready}), 
		.data_out_bus({start_0_out1_data}), .valid_out_bus({start_0_out1_valid}), .ready_out_bus({start_0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_24
		(.clk(forkC_24_clk), .rst(forkC_24_rst),
		.data_in_bus({forkC_24_in1_data}), .valid_in_bus({forkC_24_in1_valid}), .ready_in_bus({forkC_24_in1_ready}), 
		.data_out_bus({forkC_24_out3_data, forkC_24_out2_data, forkC_24_out1_data}), .valid_out_bus({forkC_24_out3_valid, forkC_24_out2_valid, forkC_24_out1_valid}), .ready_out_bus({forkC_24_out3_ready, forkC_24_out2_ready, forkC_24_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_26
		(.clk(branchC_26_clk), .rst(branchC_26_rst),
		.data_in_bus({{branchC_26_in2_data}, branchC_26_in1_data}), .valid_in_bus({branchC_26_in2_valid, branchC_26_in1_valid}), .ready_in_bus({branchC_26_in2_ready, branchC_26_in1_ready}), 
		.data_out_bus({branchC_26_out2_data, branchC_26_out1_data}), .valid_out_bus({branchC_26_out2_valid, branchC_26_out1_valid}), .ready_out_bus({branchC_26_out2_ready, branchC_26_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_25
		(.clk(fork_25_clk), .rst(fork_25_rst),
		.data_in_bus({fork_25_in1_data}), .valid_in_bus({fork_25_in1_valid}), .ready_in_bus({fork_25_in1_ready}), 
		.data_out_bus({fork_25_out2_data, fork_25_out1_data}), .valid_out_bus({fork_25_out2_valid, fork_25_out1_valid}), .ready_out_bus({fork_25_out2_ready, fork_25_out1_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(6), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_filter
		(.clk(MC_filter_clk), .rst(MC_filter_rst),
		.io_storeDataOut(filter_dout0), .io_storeAddrOut(filter_address0), .io_storeEnable(filter_we0),
		.io_loadDataIn(filter_din1), .io_loadAddrOut(filter_address1), .io_loadEnable(filter_ce1),
		.io_bbpValids({MC_filter_in2_valid}), .io_bb_stCountArray({MC_filter_in2_data}), .io_bbReadyToPrevs({MC_filter_in2_ready}), .io_rdPortsPrev_ready({MC_filter_in1_ready}), .io_rdPortsPrev_valid({MC_filter_in1_valid}), .io_rdPortsPrev_bits({MC_filter_in1_data}), 	
	.io_wrAddrPorts_ready({MC_filter_in3_ready}), .io_wrAddrPorts_valid({MC_filter_in3_valid}), .io_wrAddrPorts_bits({MC_filter_in3_data}), 	
	.io_wrDataPorts_ready({MC_filter_in4_ready}), .io_wrDataPorts_valid({MC_filter_in4_valid}), .io_wrDataPorts_bits({MC_filter_in4_data}), 	
	.io_rdPortsNext_ready({MC_filter_out1_ready}), .io_rdPortsNext_valid({MC_filter_out1_valid}), .io_rdPortsNext_bits({MC_filter_out1_data}), 	
	.io_Empty_Valid({MC_filter_out2_valid}), .io_Empty_Ready({MC_filter_out2_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(13), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_orig
		(.clk(MC_orig_clk), .rst(MC_orig_rst),
		.io_storeDataOut(orig_dout0), .io_storeAddrOut(orig_address0), .io_storeEnable(orig_we0),
		.io_loadDataIn(orig_din1), .io_loadAddrOut(orig_address1), .io_loadEnable(orig_ce1),
		.io_bbpValids({MC_orig_in2_valid}), .io_bb_stCountArray({MC_orig_in2_data}), .io_bbReadyToPrevs({MC_orig_in2_ready}), .io_rdPortsPrev_ready({MC_orig_in1_ready}), .io_rdPortsPrev_valid({MC_orig_in1_valid}), .io_rdPortsPrev_bits({MC_orig_in1_data}), 	
	.io_wrAddrPorts_ready({MC_orig_in3_ready}), .io_wrAddrPorts_valid({MC_orig_in3_valid}), .io_wrAddrPorts_bits({MC_orig_in3_data}), 	
	.io_wrDataPorts_ready({MC_orig_in4_ready}), .io_wrDataPorts_valid({MC_orig_in4_valid}), .io_wrDataPorts_bits({MC_orig_in4_data}), 	
	.io_rdPortsNext_ready({MC_orig_out1_ready}), .io_rdPortsNext_valid({MC_orig_out1_valid}), .io_rdPortsNext_bits({MC_orig_out1_data}), 	
	.io_Empty_Valid({MC_orig_out2_valid}), .io_Empty_Ready({MC_orig_out2_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(11), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_sol
		(.clk(MC_sol_clk), .rst(MC_sol_rst),
		.io_storeDataOut(sol_dout0), .io_storeAddrOut(sol_address0), .io_storeEnable(sol_we0),
		.io_loadDataIn(sol_din1), .io_loadAddrOut(sol_address1), .io_loadEnable(sol_ce1),
		.io_bbpValids({MC_sol_in1_valid}), .io_bb_stCountArray({MC_sol_in1_data}), .io_bbReadyToPrevs({MC_sol_in1_ready}), .io_rdPortsPrev_ready({MC_sol_in4_ready}), .io_rdPortsPrev_valid({MC_sol_in4_valid}), .io_rdPortsPrev_bits({MC_sol_in4_data}), 	
	.io_wrAddrPorts_ready({MC_sol_in2_ready}), .io_wrAddrPorts_valid({MC_sol_in2_valid}), .io_wrAddrPorts_bits({MC_sol_in2_data}), 	
	.io_wrDataPorts_ready({MC_sol_in3_ready}), .io_wrDataPorts_valid({MC_sol_in3_valid}), .io_wrDataPorts_bits({MC_sol_in3_data}), 	
	.io_rdPortsNext_ready({MC_sol_out2_ready}), .io_rdPortsNext_valid({MC_sol_out2_valid}), .io_rdPortsNext_bits({MC_sol_out2_data}), 	
	.io_Empty_Valid({MC_sol_out1_valid}), .io_Empty_Ready({MC_sol_out1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_1
		(.clk(sink_1_clk), .rst(sink_1_rst),
		.data_in_bus({sink_1_in1_data}), .valid_in_bus({sink_1_in1_valid}), .ready_in_bus({sink_1_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_2
		(.clk(sink_2_clk), .rst(sink_2_rst),
		.data_in_bus({sink_2_in1_data}), .valid_in_bus({sink_2_in1_valid}), .ready_in_bus({sink_2_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_3
		(.clk(sink_3_clk), .rst(sink_3_rst),
		.data_in_bus({sink_3_in1_data}), .valid_in_bus({sink_3_in1_valid}), .ready_in_bus({sink_3_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_4
		(.clk(sink_4_clk), .rst(sink_4_rst),
		.data_in_bus({sink_4_in1_data}), .valid_in_bus({sink_4_in1_valid}), .ready_in_bus({sink_4_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_5
		(.clk(sink_5_clk), .rst(sink_5_rst),
		.data_in_bus({sink_5_in1_data}), .valid_in_bus({sink_5_in1_valid}), .ready_in_bus({sink_5_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_6
		(.clk(sink_6_clk), .rst(sink_6_rst),
		.data_in_bus({sink_6_in1_data}), .valid_in_bus({sink_6_in1_valid}), .ready_in_bus({sink_6_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_7
		(.clk(sink_7_clk), .rst(sink_7_rst),
		.data_in_bus({sink_7_in1_data}), .valid_in_bus({sink_7_in1_valid}), .ready_in_bus({sink_7_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_8
		(.clk(sink_8_clk), .rst(sink_8_rst),
		.data_in_bus({sink_8_in1_data}), .valid_in_bus({sink_8_in1_valid}), .ready_in_bus({sink_8_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_9
		(.clk(sink_9_clk), .rst(sink_9_rst),
		.data_in_bus({sink_9_in1_data}), .valid_in_bus({sink_9_in1_valid}), .ready_in_bus({sink_9_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(3))sink_node_sink_10
		(.clk(sink_10_clk), .rst(sink_10_rst),
		.data_in_bus({sink_10_in1_data}), .valid_in_bus({sink_10_in1_valid}), .ready_in_bus({sink_10_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_11
		(.clk(sink_11_clk), .rst(sink_11_rst),
		.data_in_bus({sink_11_in1_data}), .valid_in_bus({sink_11_in1_valid}), .ready_in_bus({sink_11_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_12
		(.clk(sink_12_clk), .rst(sink_12_rst),
		.data_in_bus({sink_12_in1_data}), .valid_in_bus({sink_12_in1_valid}), .ready_in_bus({sink_12_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(3))sink_node_sink_13
		(.clk(sink_13_clk), .rst(sink_13_rst),
		.data_in_bus({sink_13_in1_data}), .valid_in_bus({sink_13_in1_valid}), .ready_in_bus({sink_13_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(3))sink_node_sink_14
		(.clk(sink_14_clk), .rst(sink_14_rst),
		.data_in_bus({sink_14_in1_data}), .valid_in_bus({sink_14_in1_valid}), .ready_in_bus({sink_14_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_15
		(.clk(sink_15_clk), .rst(sink_15_rst),
		.data_in_bus({sink_15_in1_data}), .valid_in_bus({sink_15_in1_valid}), .ready_in_bus({sink_15_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_16
		(.clk(sink_16_clk), .rst(sink_16_rst),
		.data_in_bus({sink_16_in1_data}), .valid_in_bus({sink_16_in1_valid}), .ready_in_bus({sink_16_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_17
		(.clk(sink_17_clk), .rst(sink_17_rst),
		.data_in_bus({sink_17_in1_data}), .valid_in_bus({sink_17_in1_valid}), .ready_in_bus({sink_17_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(5))sink_node_sink_18
		(.clk(sink_18_clk), .rst(sink_18_rst),
		.data_in_bus({sink_18_in1_data}), .valid_in_bus({sink_18_in1_valid}), .ready_in_bus({sink_18_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_19
		(.clk(sink_19_clk), .rst(sink_19_rst),
		.data_in_bus({sink_19_in1_data}), .valid_in_bus({sink_19_in1_valid}), .ready_in_bus({sink_19_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_20
		(.clk(sink_20_clk), .rst(sink_20_rst),
		.data_in_bus({sink_20_in1_data}), .valid_in_bus({sink_20_in1_valid}), .ready_in_bus({sink_20_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_21
		(.clk(sink_21_clk), .rst(sink_21_rst),
		.data_in_bus({sink_21_in1_data}), .valid_in_bus({sink_21_in1_valid}), .ready_in_bus({sink_21_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_22
		(.clk(sink_22_clk), .rst(sink_22_rst),
		.data_in_bus({sink_22_in1_data}), .valid_in_bus({sink_22_in1_valid}), .ready_in_bus({sink_22_in1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_100
		(.clk(Buffer_100_clk), .rst(Buffer_100_rst),
		.data_in_bus({Buffer_100_in1_data}), .valid_in_bus({Buffer_100_in1_valid}), .ready_in_bus({Buffer_100_in1_ready}), 
		.data_out_bus({Buffer_100_out1_data}), .valid_out_bus({Buffer_100_out1_valid}), .ready_out_bus({Buffer_100_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_101
		(.clk(Buffer_101_clk), .rst(Buffer_101_rst),
		.data_in_bus({Buffer_101_in1_data}), .valid_in_bus({Buffer_101_in1_valid}), .ready_in_bus({Buffer_101_in1_ready}), 
		.data_out_bus({Buffer_101_out1_data}), .valid_out_bus({Buffer_101_out1_valid}), .ready_out_bus({Buffer_101_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_102
		(.clk(Buffer_102_clk), .rst(Buffer_102_rst),
		.data_in_bus({Buffer_102_in1_data}), .valid_in_bus({Buffer_102_in1_valid}), .ready_in_bus({Buffer_102_in1_ready}), 
		.data_out_bus({Buffer_102_out1_data}), .valid_out_bus({Buffer_102_out1_valid}), .ready_out_bus({Buffer_102_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_103
		(.clk(Buffer_103_clk), .rst(Buffer_103_rst),
		.data_in_bus({Buffer_103_in1_data}), .valid_in_bus({Buffer_103_in1_valid}), .ready_in_bus({Buffer_103_in1_ready}), 
		.data_out_bus({Buffer_103_out1_data}), .valid_out_bus({Buffer_103_out1_valid}), .ready_out_bus({Buffer_103_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_104
		(.clk(Buffer_104_clk), .rst(Buffer_104_rst),
		.data_in_bus({Buffer_104_in1_data}), .valid_in_bus({Buffer_104_in1_valid}), .ready_in_bus({Buffer_104_in1_ready}), 
		.data_out_bus({Buffer_104_out1_data}), .valid_out_bus({Buffer_104_out1_valid}), .ready_out_bus({Buffer_104_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_105
		(.clk(Buffer_105_clk), .rst(Buffer_105_rst),
		.data_in_bus({Buffer_105_in1_data}), .valid_in_bus({Buffer_105_in1_valid}), .ready_in_bus({Buffer_105_in1_ready}), 
		.data_out_bus({Buffer_105_out1_data}), .valid_out_bus({Buffer_105_out1_valid}), .ready_out_bus({Buffer_105_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_106
		(.clk(Buffer_106_clk), .rst(Buffer_106_rst),
		.data_in_bus({Buffer_106_in1_data}), .valid_in_bus({Buffer_106_in1_valid}), .ready_in_bus({Buffer_106_in1_ready}), 
		.data_out_bus({Buffer_106_out1_data}), .valid_out_bus({Buffer_106_out1_valid}), .ready_out_bus({Buffer_106_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_107
		(.clk(Buffer_107_clk), .rst(Buffer_107_rst),
		.data_in_bus({Buffer_107_in1_data}), .valid_in_bus({Buffer_107_in1_valid}), .ready_in_bus({Buffer_107_in1_ready}), 
		.data_out_bus({Buffer_107_out1_data}), .valid_out_bus({Buffer_107_out1_valid}), .ready_out_bus({Buffer_107_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_108
		(.clk(Buffer_108_clk), .rst(Buffer_108_rst),
		.data_in_bus({Buffer_108_in1_data}), .valid_in_bus({Buffer_108_in1_valid}), .ready_in_bus({Buffer_108_in1_ready}), 
		.data_out_bus({Buffer_108_out1_data}), .valid_out_bus({Buffer_108_out1_valid}), .ready_out_bus({Buffer_108_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_109
		(.clk(Buffer_109_clk), .rst(Buffer_109_rst),
		.data_in_bus({Buffer_109_in1_data}), .valid_in_bus({Buffer_109_in1_valid}), .ready_in_bus({Buffer_109_in1_ready}), 
		.data_out_bus({Buffer_109_out1_data}), .valid_out_bus({Buffer_109_out1_valid}), .ready_out_bus({Buffer_109_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_110
		(.clk(Buffer_110_clk), .rst(Buffer_110_rst),
		.data_in_bus({Buffer_110_in1_data}), .valid_in_bus({Buffer_110_in1_valid}), .ready_in_bus({Buffer_110_in1_ready}), 
		.data_out_bus({Buffer_110_out1_data}), .valid_out_bus({Buffer_110_out1_valid}), .ready_out_bus({Buffer_110_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_111
		(.clk(Buffer_111_clk), .rst(Buffer_111_rst),
		.data_in_bus({Buffer_111_in1_data}), .valid_in_bus({Buffer_111_in1_valid}), .ready_in_bus({Buffer_111_in1_ready}), 
		.data_out_bus({Buffer_111_out1_data}), .valid_out_bus({Buffer_111_out1_valid}), .ready_out_bus({Buffer_111_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_112
		(.clk(Buffer_112_clk), .rst(Buffer_112_rst),
		.data_in_bus({Buffer_112_in1_data}), .valid_in_bus({Buffer_112_in1_valid}), .ready_in_bus({Buffer_112_in1_ready}), 
		.data_out_bus({Buffer_112_out1_data}), .valid_out_bus({Buffer_112_out1_valid}), .ready_out_bus({Buffer_112_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_113
		(.clk(Buffer_113_clk), .rst(Buffer_113_rst),
		.data_in_bus({Buffer_113_in1_data}), .valid_in_bus({Buffer_113_in1_valid}), .ready_in_bus({Buffer_113_in1_ready}), 
		.data_out_bus({Buffer_113_out1_data}), .valid_out_bus({Buffer_113_out1_valid}), .ready_out_bus({Buffer_113_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_114
		(.clk(Buffer_114_clk), .rst(Buffer_114_rst),
		.data_in_bus({Buffer_114_in1_data}), .valid_in_bus({Buffer_114_in1_valid}), .ready_in_bus({Buffer_114_in1_ready}), 
		.data_out_bus({Buffer_114_out1_data}), .valid_out_bus({Buffer_114_out1_valid}), .ready_out_bus({Buffer_114_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_115
		(.clk(Buffer_115_clk), .rst(Buffer_115_rst),
		.data_in_bus({Buffer_115_in1_data}), .valid_in_bus({Buffer_115_in1_valid}), .ready_in_bus({Buffer_115_in1_ready}), 
		.data_out_bus({Buffer_115_out1_data}), .valid_out_bus({Buffer_115_out1_valid}), .ready_out_bus({Buffer_115_out1_ready}));

endmodule

