module matrix(
	input clk,
	input rst,

	input [0 : 0]start_in,
	input start_valid,
	output start_ready,

	output [0 : 0]end_out,
	output end_valid,
	input end_ready,

	output [11 : 0]in_a_address0,
	output in_a_ce0,
	output in_a_we0,
	output [31 : 0]in_a_dout0,
	input [31 : 0]in_a_din0,
	output [11 : 0]in_a_address1,
	output in_a_ce1,
	output in_a_we1,
	output [31 : 0]in_a_dout1,
	input [31 : 0]in_a_din1,

	output [11 : 0]in_b_address0,
	output in_b_ce0,
	output in_b_we0,
	output [31 : 0]in_b_dout0,
	input [31 : 0]in_b_din0,
	output [11 : 0]in_b_address1,
	output in_b_ce1,
	output in_b_we1,
	output [31 : 0]in_b_dout1,
	input [31 : 0]in_b_din1,

	output [11 : 0]out_c_address0,
	output out_c_ce0,
	output out_c_we0,
	output [31 : 0]out_c_dout0,
	input [31 : 0]out_c_din0,
	output [11 : 0]out_c_address1,
	output out_c_ce1,
	output out_c_we1,
	output [31 : 0]out_c_dout1,
	input [31 : 0]out_c_din1

);

	wire brCst_block1_clk;
	wire brCst_block1_rst;
	wire [0 : 0]brCst_block1_in1_data;
	wire brCst_block1_in1_ready;
	wire brCst_block1_in1_valid;
	wire [0 : 0]brCst_block1_out1_data;
	wire brCst_block1_out1_ready;
	wire brCst_block1_out1_valid;

	wire cst_0_clk;
	wire cst_0_rst;
	wire [0 : 0]cst_0_in1_data;
	wire cst_0_in1_ready;
	wire cst_0_in1_valid;
	wire [0 : 0]cst_0_out1_data;
	wire cst_0_out1_ready;
	wire cst_0_out1_valid;

	wire branch_0_clk;
	wire branch_0_rst;
	wire [0 : 0]branch_0_in1_data;
	wire branch_0_in1_ready;
	wire branch_0_in1_valid;
	wire [0 : 0]branch_0_in2_data;
	wire branch_0_in2_ready;
	wire branch_0_in2_valid;
	wire [0 : 0]branch_0_out1_data;
	wire branch_0_out1_ready;
	wire branch_0_out1_valid;
	wire [0 : 0]branch_0_out2_data;
	wire branch_0_out2_ready;
	wire branch_0_out2_valid;

	wire start_0_clk;
	wire start_0_rst;
	wire [0 : 0]start_0_in1_data;
	wire start_0_in1_ready;
	wire start_0_in1_valid;
	wire [0 : 0]start_0_out1_data;
	wire start_0_out1_ready;
	wire start_0_out1_valid;

	wire forkC_16_clk;
	wire forkC_16_rst;
	wire [0 : 0]forkC_16_in1_data;
	wire forkC_16_in1_ready;
	wire forkC_16_in1_valid;
	wire [0 : 0]forkC_16_out1_data;
	wire forkC_16_out1_ready;
	wire forkC_16_out1_valid;
	wire [0 : 0]forkC_16_out2_data;
	wire forkC_16_out2_ready;
	wire forkC_16_out2_valid;
	wire [0 : 0]forkC_16_out3_data;
	wire forkC_16_out3_ready;
	wire forkC_16_out3_valid;

	wire branchC_14_clk;
	wire branchC_14_rst;
	wire [0 : 0]branchC_14_in1_data;
	wire branchC_14_in1_ready;
	wire branchC_14_in1_valid;
	wire [0 : 0]branchC_14_in2_data;
	wire branchC_14_in2_ready;
	wire branchC_14_in2_valid;
	wire [0 : 0]branchC_14_out1_data;
	wire branchC_14_out1_ready;
	wire branchC_14_out1_valid;
	wire [0 : 0]branchC_14_out2_data;
	wire branchC_14_out2_ready;
	wire branchC_14_out2_valid;

	wire fork_17_clk;
	wire fork_17_rst;
	wire [0 : 0]fork_17_in1_data;
	wire fork_17_in1_ready;
	wire fork_17_in1_valid;
	wire [0 : 0]fork_17_out1_data;
	wire fork_17_out1_ready;
	wire fork_17_out1_valid;
	wire [0 : 0]fork_17_out2_data;
	wire fork_17_out2_ready;
	wire fork_17_out2_valid;

	wire phi_3_clk;
	wire phi_3_rst;
	wire [0 : 0]phi_3_in1_data;
	wire phi_3_in1_ready;
	wire phi_3_in1_valid;
	wire [5 : 0]phi_3_in2_data;
	wire phi_3_in2_ready;
	wire phi_3_in2_valid;
	wire [5 : 0]phi_3_in3_data;
	wire phi_3_in3_ready;
	wire phi_3_in3_valid;
	wire [5 : 0]phi_3_out1_data;
	wire phi_3_out1_ready;
	wire phi_3_out1_valid;

	wire brCst_block3_clk;
	wire brCst_block3_rst;
	wire [0 : 0]brCst_block3_in1_data;
	wire brCst_block3_in1_ready;
	wire brCst_block3_in1_valid;
	wire [0 : 0]brCst_block3_out1_data;
	wire brCst_block3_out1_ready;
	wire brCst_block3_out1_valid;

	wire cst_2_clk;
	wire cst_2_rst;
	wire [0 : 0]cst_2_in1_data;
	wire cst_2_in1_ready;
	wire cst_2_in1_valid;
	wire [0 : 0]cst_2_out1_data;
	wire cst_2_out1_ready;
	wire cst_2_out1_valid;

	wire cst_3_clk;
	wire cst_3_rst;
	wire [0 : 0]cst_3_in1_data;
	wire cst_3_in1_ready;
	wire cst_3_in1_valid;
	wire [0 : 0]cst_3_out1_data;
	wire cst_3_out1_ready;
	wire cst_3_out1_valid;

	wire phi_n1_clk;
	wire phi_n1_rst;
	wire [5 : 0]phi_n1_in1_data;
	wire phi_n1_in1_ready;
	wire phi_n1_in1_valid;
	wire [5 : 0]phi_n1_in2_data;
	wire phi_n1_in2_ready;
	wire phi_n1_in2_valid;
	wire [5 : 0]phi_n1_out1_data;
	wire phi_n1_out1_ready;
	wire phi_n1_out1_valid;

	wire branch_3_clk;
	wire branch_3_rst;
	wire [0 : 0]branch_3_in1_data;
	wire branch_3_in1_ready;
	wire branch_3_in1_valid;
	wire [0 : 0]branch_3_in2_data;
	wire branch_3_in2_ready;
	wire branch_3_in2_valid;
	wire [0 : 0]branch_3_out1_data;
	wire branch_3_out1_ready;
	wire branch_3_out1_valid;
	wire [0 : 0]branch_3_out2_data;
	wire branch_3_out2_ready;
	wire branch_3_out2_valid;

	wire branch_4_clk;
	wire branch_4_rst;
	wire [0 : 0]branch_4_in1_data;
	wire branch_4_in1_ready;
	wire branch_4_in1_valid;
	wire [0 : 0]branch_4_in2_data;
	wire branch_4_in2_ready;
	wire branch_4_in2_valid;
	wire [0 : 0]branch_4_out1_data;
	wire branch_4_out1_ready;
	wire branch_4_out1_valid;
	wire [0 : 0]branch_4_out2_data;
	wire branch_4_out2_ready;
	wire branch_4_out2_valid;

	wire branch_5_clk;
	wire branch_5_rst;
	wire [5 : 0]branch_5_in1_data;
	wire branch_5_in1_ready;
	wire branch_5_in1_valid;
	wire [0 : 0]branch_5_in2_data;
	wire branch_5_in2_ready;
	wire branch_5_in2_valid;
	wire [5 : 0]branch_5_out1_data;
	wire branch_5_out1_ready;
	wire branch_5_out1_valid;
	wire [5 : 0]branch_5_out2_data;
	wire branch_5_out2_ready;
	wire branch_5_out2_valid;

	wire branch_6_clk;
	wire branch_6_rst;
	wire [5 : 0]branch_6_in1_data;
	wire branch_6_in1_ready;
	wire branch_6_in1_valid;
	wire [0 : 0]branch_6_in2_data;
	wire branch_6_in2_ready;
	wire branch_6_in2_valid;
	wire [5 : 0]branch_6_out1_data;
	wire branch_6_out1_ready;
	wire branch_6_out1_valid;
	wire [5 : 0]branch_6_out2_data;
	wire branch_6_out2_ready;
	wire branch_6_out2_valid;

	wire fork_11_clk;
	wire fork_11_rst;
	wire [0 : 0]fork_11_in1_data;
	wire fork_11_in1_ready;
	wire fork_11_in1_valid;
	wire [0 : 0]fork_11_out1_data;
	wire fork_11_out1_ready;
	wire fork_11_out1_valid;
	wire [0 : 0]fork_11_out2_data;
	wire fork_11_out2_ready;
	wire fork_11_out2_valid;
	wire [0 : 0]fork_11_out3_data;
	wire fork_11_out3_ready;
	wire fork_11_out3_valid;
	wire [0 : 0]fork_11_out4_data;
	wire fork_11_out4_ready;
	wire fork_11_out4_valid;
	wire [0 : 0]fork_11_out5_data;
	wire fork_11_out5_ready;
	wire fork_11_out5_valid;

	wire phiC_8_clk;
	wire phiC_8_rst;
	wire [0 : 0]phiC_8_in1_data;
	wire phiC_8_in1_ready;
	wire phiC_8_in1_valid;
	wire [0 : 0]phiC_8_in2_data;
	wire phiC_8_in2_ready;
	wire phiC_8_in2_valid;
	wire [0 : 0]phiC_8_out1_data;
	wire phiC_8_out1_ready;
	wire phiC_8_out1_valid;
	wire [0 : 0]phiC_8_out2_data;
	wire phiC_8_out2_ready;
	wire phiC_8_out2_valid;

	wire forkC_19_clk;
	wire forkC_19_rst;
	wire [0 : 0]forkC_19_in1_data;
	wire forkC_19_in1_ready;
	wire forkC_19_in1_valid;
	wire [0 : 0]forkC_19_out1_data;
	wire forkC_19_out1_ready;
	wire forkC_19_out1_valid;
	wire [0 : 0]forkC_19_out2_data;
	wire forkC_19_out2_ready;
	wire forkC_19_out2_valid;
	wire [0 : 0]forkC_19_out3_data;
	wire forkC_19_out3_ready;
	wire forkC_19_out3_valid;
	wire [0 : 0]forkC_19_out4_data;
	wire forkC_19_out4_ready;
	wire forkC_19_out4_valid;

	wire branchC_16_clk;
	wire branchC_16_rst;
	wire [0 : 0]branchC_16_in1_data;
	wire branchC_16_in1_ready;
	wire branchC_16_in1_valid;
	wire [0 : 0]branchC_16_in2_data;
	wire branchC_16_in2_ready;
	wire branchC_16_in2_valid;
	wire [0 : 0]branchC_16_out1_data;
	wire branchC_16_out1_ready;
	wire branchC_16_out1_valid;
	wire [0 : 0]branchC_16_out2_data;
	wire branchC_16_out2_ready;
	wire branchC_16_out2_valid;

	wire cst_11_clk;
	wire cst_11_rst;
	wire [0 : 0]cst_11_in1_data;
	wire cst_11_in1_ready;
	wire cst_11_in1_valid;
	wire [0 : 0]cst_11_out1_data;
	wire cst_11_out1_ready;
	wire cst_11_out1_valid;

	wire add_29_clk;
	wire add_29_rst;
	wire [5 : 0]add_29_in1_data;
	wire add_29_in1_ready;
	wire add_29_in1_valid;
	wire [5 : 0]add_29_in2_data;
	wire add_29_in2_ready;
	wire add_29_in2_valid;
	wire [5 : 0]add_29_out1_data;
	wire add_29_out1_ready;
	wire add_29_out1_valid;

	wire cst_12_clk;
	wire cst_12_rst;
	wire [5 : 0]cst_12_in1_data;
	wire cst_12_in1_ready;
	wire cst_12_in1_valid;
	wire [5 : 0]cst_12_out1_data;
	wire cst_12_out1_ready;
	wire cst_12_out1_valid;

	wire icmp_30_clk;
	wire icmp_30_rst;
	wire [5 : 0]icmp_30_in1_data;
	wire icmp_30_in1_ready;
	wire icmp_30_in1_valid;
	wire [5 : 0]icmp_30_in2_data;
	wire icmp_30_in2_ready;
	wire icmp_30_in2_valid;
	wire [0 : 0]icmp_30_out1_data;
	wire icmp_30_out1_ready;
	wire icmp_30_out1_valid;

	wire phi_n0_clk;
	wire phi_n0_rst;
	wire [5 : 0]phi_n0_in1_data;
	wire phi_n0_in1_ready;
	wire phi_n0_in1_valid;
	wire [5 : 0]phi_n0_out1_data;
	wire phi_n0_out1_ready;
	wire phi_n0_out1_valid;

	wire fork_4_clk;
	wire fork_4_rst;
	wire [5 : 0]fork_4_in1_data;
	wire fork_4_in1_ready;
	wire fork_4_in1_valid;
	wire [5 : 0]fork_4_out1_data;
	wire fork_4_out1_ready;
	wire fork_4_out1_valid;
	wire [5 : 0]fork_4_out2_data;
	wire fork_4_out2_ready;
	wire fork_4_out2_valid;

	wire branch_13_clk;
	wire branch_13_rst;
	wire [5 : 0]branch_13_in1_data;
	wire branch_13_in1_ready;
	wire branch_13_in1_valid;
	wire [0 : 0]branch_13_in2_data;
	wire branch_13_in2_ready;
	wire branch_13_in2_valid;
	wire [5 : 0]branch_13_out1_data;
	wire branch_13_out1_ready;
	wire branch_13_out1_valid;
	wire [5 : 0]branch_13_out2_data;
	wire branch_13_out2_ready;
	wire branch_13_out2_valid;

	wire phiC_11_clk;
	wire phiC_11_rst;
	wire [0 : 0]phiC_11_in1_data;
	wire phiC_11_in1_ready;
	wire phiC_11_in1_valid;
	wire [0 : 0]phiC_11_out1_data;
	wire phiC_11_out1_ready;
	wire phiC_11_out1_valid;

	wire branchC_19_clk;
	wire branchC_19_rst;
	wire [0 : 0]branchC_19_in1_data;
	wire branchC_19_in1_ready;
	wire branchC_19_in1_valid;
	wire [0 : 0]branchC_19_in2_data;
	wire branchC_19_in2_ready;
	wire branchC_19_in2_valid;
	wire [0 : 0]branchC_19_out1_data;
	wire branchC_19_out1_ready;
	wire branchC_19_out1_valid;
	wire [0 : 0]branchC_19_out2_data;
	wire branchC_19_out2_ready;
	wire branchC_19_out2_valid;

	wire fork_23_clk;
	wire fork_23_rst;
	wire [0 : 0]fork_23_in1_data;
	wire fork_23_in1_ready;
	wire fork_23_in1_valid;
	wire [0 : 0]fork_23_out1_data;
	wire fork_23_out1_ready;
	wire fork_23_out1_valid;
	wire [0 : 0]fork_23_out2_data;
	wire fork_23_out2_ready;
	wire fork_23_out2_valid;

	wire source_7_clk;
	wire source_7_rst;
	wire [0 : 0]source_7_out1_data;
	wire source_7_out1_ready;
	wire source_7_out1_valid;

	wire source_8_clk;
	wire source_8_rst;
	wire [5 : 0]source_8_out1_data;
	wire source_8_out1_ready;
	wire source_8_out1_valid;

	wire phi_5_clk;
	wire phi_5_rst;
	wire [0 : 0]phi_5_in1_data;
	wire phi_5_in1_ready;
	wire phi_5_in1_valid;
	wire [31 : 0]phi_5_in2_data;
	wire phi_5_in2_ready;
	wire phi_5_in2_valid;
	wire [31 : 0]phi_5_in3_data;
	wire phi_5_in3_ready;
	wire phi_5_in3_valid;
	wire [31 : 0]phi_5_out1_data;
	wire phi_5_out1_ready;
	wire phi_5_out1_valid;

	wire phi_6_clk;
	wire phi_6_rst;
	wire [0 : 0]phi_6_in1_data;
	wire phi_6_in1_ready;
	wire phi_6_in1_valid;
	wire [5 : 0]phi_6_in2_data;
	wire phi_6_in2_ready;
	wire phi_6_in2_valid;
	wire [5 : 0]phi_6_in3_data;
	wire phi_6_in3_ready;
	wire phi_6_in3_valid;
	wire [5 : 0]phi_6_out1_data;
	wire phi_6_out1_ready;
	wire phi_6_out1_valid;

	wire cst_4_clk;
	wire cst_4_rst;
	wire [2 : 0]cst_4_in1_data;
	wire cst_4_in1_ready;
	wire cst_4_in1_valid;
	wire [2 : 0]cst_4_out1_data;
	wire cst_4_out1_ready;
	wire cst_4_out1_valid;

	wire shl_7_clk;
	wire shl_7_rst;
	wire [10 : 0]shl_7_in1_data;
	wire shl_7_in1_ready;
	wire shl_7_in1_valid;
	wire [10 : 0]shl_7_in2_data;
	wire shl_7_in2_ready;
	wire shl_7_in2_valid;
	wire [10 : 0]shl_7_out1_data;
	wire shl_7_out1_ready;
	wire shl_7_out1_valid;

	wire add_8_clk;
	wire add_8_rst;
	wire [11 : 0]add_8_in1_data;
	wire add_8_in1_ready;
	wire add_8_in1_valid;
	wire [11 : 0]add_8_in2_data;
	wire add_8_in2_ready;
	wire add_8_in2_valid;
	wire [11 : 0]add_8_out1_data;
	wire add_8_out1_ready;
	wire add_8_out1_valid;

	wire load_11_clk;
	wire load_11_rst;
	wire [31 : 0]load_11_in1_data;
	wire load_11_in1_ready;
	wire load_11_in1_valid;
	wire [11 : 0]load_11_in2_data;
	wire load_11_in2_ready;
	wire load_11_in2_valid;
	wire [31 : 0]load_11_out1_data;
	wire load_11_out1_ready;
	wire load_11_out1_valid;
	wire [11 : 0]load_11_out2_data;
	wire load_11_out2_ready;
	wire load_11_out2_valid;

	wire cst_5_clk;
	wire cst_5_rst;
	wire [2 : 0]cst_5_in1_data;
	wire cst_5_in1_ready;
	wire cst_5_in1_valid;
	wire [2 : 0]cst_5_out1_data;
	wire cst_5_out1_ready;
	wire cst_5_out1_valid;

	wire shl_12_clk;
	wire shl_12_rst;
	wire [10 : 0]shl_12_in1_data;
	wire shl_12_in1_ready;
	wire shl_12_in1_valid;
	wire [10 : 0]shl_12_in2_data;
	wire shl_12_in2_ready;
	wire shl_12_in2_valid;
	wire [10 : 0]shl_12_out1_data;
	wire shl_12_out1_ready;
	wire shl_12_out1_valid;

	wire add_13_clk;
	wire add_13_rst;
	wire [11 : 0]add_13_in1_data;
	wire add_13_in1_ready;
	wire add_13_in1_valid;
	wire [11 : 0]add_13_in2_data;
	wire add_13_in2_ready;
	wire add_13_in2_valid;
	wire [11 : 0]add_13_out1_data;
	wire add_13_out1_ready;
	wire add_13_out1_valid;

	wire load_16_clk;
	wire load_16_rst;
	wire [31 : 0]load_16_in1_data;
	wire load_16_in1_ready;
	wire load_16_in1_valid;
	wire [11 : 0]load_16_in2_data;
	wire load_16_in2_ready;
	wire load_16_in2_valid;
	wire [31 : 0]load_16_out1_data;
	wire load_16_out1_ready;
	wire load_16_out1_valid;
	wire [11 : 0]load_16_out2_data;
	wire load_16_out2_ready;
	wire load_16_out2_valid;

	wire mul_17_clk;
	wire mul_17_rst;
	wire [15 : 0]mul_17_in1_data;
	wire mul_17_in1_ready;
	wire mul_17_in1_valid;
	wire [15 : 0]mul_17_in2_data;
	wire mul_17_in2_ready;
	wire mul_17_in2_valid;
	wire [31 : 0]mul_17_out1_data;
	wire mul_17_out1_ready;
	wire mul_17_out1_valid;

	wire add_18_clk;
	wire add_18_rst;
	wire [31 : 0]add_18_in1_data;
	wire add_18_in1_ready;
	wire add_18_in1_valid;
	wire [31 : 0]add_18_in2_data;
	wire add_18_in2_ready;
	wire add_18_in2_valid;
	wire [31 : 0]add_18_out1_data;
	wire add_18_out1_ready;
	wire add_18_out1_valid;

	wire cst_6_clk;
	wire cst_6_rst;
	wire [0 : 0]cst_6_in1_data;
	wire cst_6_in1_ready;
	wire cst_6_in1_valid;
	wire [0 : 0]cst_6_out1_data;
	wire cst_6_out1_ready;
	wire cst_6_out1_valid;

	wire add_19_clk;
	wire add_19_rst;
	wire [5 : 0]add_19_in1_data;
	wire add_19_in1_ready;
	wire add_19_in1_valid;
	wire [5 : 0]add_19_in2_data;
	wire add_19_in2_ready;
	wire add_19_in2_valid;
	wire [5 : 0]add_19_out1_data;
	wire add_19_out1_ready;
	wire add_19_out1_valid;

	wire cst_7_clk;
	wire cst_7_rst;
	wire [5 : 0]cst_7_in1_data;
	wire cst_7_in1_ready;
	wire cst_7_in1_valid;
	wire [5 : 0]cst_7_out1_data;
	wire cst_7_out1_ready;
	wire cst_7_out1_valid;

	wire icmp_20_clk;
	wire icmp_20_rst;
	wire [5 : 0]icmp_20_in1_data;
	wire icmp_20_in1_ready;
	wire icmp_20_in1_valid;
	wire [5 : 0]icmp_20_in2_data;
	wire icmp_20_in2_ready;
	wire icmp_20_in2_valid;
	wire [0 : 0]icmp_20_out1_data;
	wire icmp_20_out1_ready;
	wire icmp_20_out1_valid;

	wire phi_n5_clk;
	wire phi_n5_rst;
	wire [5 : 0]phi_n5_in1_data;
	wire phi_n5_in1_ready;
	wire phi_n5_in1_valid;
	wire [5 : 0]phi_n5_in2_data;
	wire phi_n5_in2_ready;
	wire phi_n5_in2_valid;
	wire [5 : 0]phi_n5_out1_data;
	wire phi_n5_out1_ready;
	wire phi_n5_out1_valid;

	wire phi_n6_clk;
	wire phi_n6_rst;
	wire [5 : 0]phi_n6_in1_data;
	wire phi_n6_in1_ready;
	wire phi_n6_in1_valid;
	wire [5 : 0]phi_n6_in2_data;
	wire phi_n6_in2_ready;
	wire phi_n6_in2_valid;
	wire [5 : 0]phi_n6_out1_data;
	wire phi_n6_out1_ready;
	wire phi_n6_out1_valid;

	wire fork_0_clk;
	wire fork_0_rst;
	wire [5 : 0]fork_0_in1_data;
	wire fork_0_in1_ready;
	wire fork_0_in1_valid;
	wire [5 : 0]fork_0_out1_data;
	wire fork_0_out1_ready;
	wire fork_0_out1_valid;
	wire [5 : 0]fork_0_out2_data;
	wire fork_0_out2_ready;
	wire fork_0_out2_valid;
	wire [5 : 0]fork_0_out3_data;
	wire fork_0_out3_ready;
	wire fork_0_out3_valid;

	wire fork_2_clk;
	wire fork_2_rst;
	wire [5 : 0]fork_2_in1_data;
	wire fork_2_in1_ready;
	wire fork_2_in1_valid;
	wire [5 : 0]fork_2_out1_data;
	wire fork_2_out1_ready;
	wire fork_2_out1_valid;
	wire [5 : 0]fork_2_out2_data;
	wire fork_2_out2_ready;
	wire fork_2_out2_valid;

	wire fork_7_clk;
	wire fork_7_rst;
	wire [5 : 0]fork_7_in1_data;
	wire fork_7_in1_ready;
	wire fork_7_in1_valid;
	wire [5 : 0]fork_7_out1_data;
	wire fork_7_out1_ready;
	wire fork_7_out1_valid;
	wire [5 : 0]fork_7_out2_data;
	wire fork_7_out2_ready;
	wire fork_7_out2_valid;

	wire fork_8_clk;
	wire fork_8_rst;
	wire [5 : 0]fork_8_in1_data;
	wire fork_8_in1_ready;
	wire fork_8_in1_valid;
	wire [5 : 0]fork_8_out1_data;
	wire fork_8_out1_ready;
	wire fork_8_out1_valid;
	wire [5 : 0]fork_8_out2_data;
	wire fork_8_out2_ready;
	wire fork_8_out2_valid;

	wire branch_7_clk;
	wire branch_7_rst;
	wire [31 : 0]branch_7_in1_data;
	wire branch_7_in1_ready;
	wire branch_7_in1_valid;
	wire [0 : 0]branch_7_in2_data;
	wire branch_7_in2_ready;
	wire branch_7_in2_valid;
	wire [31 : 0]branch_7_out1_data;
	wire branch_7_out1_ready;
	wire branch_7_out1_valid;
	wire [31 : 0]branch_7_out2_data;
	wire branch_7_out2_ready;
	wire branch_7_out2_valid;

	wire branch_8_clk;
	wire branch_8_rst;
	wire [5 : 0]branch_8_in1_data;
	wire branch_8_in1_ready;
	wire branch_8_in1_valid;
	wire [0 : 0]branch_8_in2_data;
	wire branch_8_in2_ready;
	wire branch_8_in2_valid;
	wire [5 : 0]branch_8_out1_data;
	wire branch_8_out1_ready;
	wire branch_8_out1_valid;
	wire [5 : 0]branch_8_out2_data;
	wire branch_8_out2_ready;
	wire branch_8_out2_valid;

	wire branch_9_clk;
	wire branch_9_rst;
	wire [5 : 0]branch_9_in1_data;
	wire branch_9_in1_ready;
	wire branch_9_in1_valid;
	wire [0 : 0]branch_9_in2_data;
	wire branch_9_in2_ready;
	wire branch_9_in2_valid;
	wire [5 : 0]branch_9_out1_data;
	wire branch_9_out1_ready;
	wire branch_9_out1_valid;
	wire [5 : 0]branch_9_out2_data;
	wire branch_9_out2_ready;
	wire branch_9_out2_valid;

	wire branch_10_clk;
	wire branch_10_rst;
	wire [5 : 0]branch_10_in1_data;
	wire branch_10_in1_ready;
	wire branch_10_in1_valid;
	wire [0 : 0]branch_10_in2_data;
	wire branch_10_in2_ready;
	wire branch_10_in2_valid;
	wire [5 : 0]branch_10_out1_data;
	wire branch_10_out1_ready;
	wire branch_10_out1_valid;
	wire [5 : 0]branch_10_out2_data;
	wire branch_10_out2_ready;
	wire branch_10_out2_valid;

	wire fork_12_clk;
	wire fork_12_rst;
	wire [0 : 0]fork_12_in1_data;
	wire fork_12_in1_ready;
	wire fork_12_in1_valid;
	wire [0 : 0]fork_12_out1_data;
	wire fork_12_out1_ready;
	wire fork_12_out1_valid;
	wire [0 : 0]fork_12_out2_data;
	wire fork_12_out2_ready;
	wire fork_12_out2_valid;
	wire [0 : 0]fork_12_out3_data;
	wire fork_12_out3_ready;
	wire fork_12_out3_valid;
	wire [0 : 0]fork_12_out4_data;
	wire fork_12_out4_ready;
	wire fork_12_out4_valid;
	wire [0 : 0]fork_12_out5_data;
	wire fork_12_out5_ready;
	wire fork_12_out5_valid;

	wire phiC_9_clk;
	wire phiC_9_rst;
	wire [0 : 0]phiC_9_in1_data;
	wire phiC_9_in1_ready;
	wire phiC_9_in1_valid;
	wire [0 : 0]phiC_9_in2_data;
	wire phiC_9_in2_ready;
	wire phiC_9_in2_valid;
	wire [0 : 0]phiC_9_out1_data;
	wire phiC_9_out1_ready;
	wire phiC_9_out1_valid;
	wire [0 : 0]phiC_9_out2_data;
	wire phiC_9_out2_ready;
	wire phiC_9_out2_valid;

	wire branchC_17_clk;
	wire branchC_17_rst;
	wire [0 : 0]branchC_17_in1_data;
	wire branchC_17_in1_ready;
	wire branchC_17_in1_valid;
	wire [0 : 0]branchC_17_in2_data;
	wire branchC_17_in2_ready;
	wire branchC_17_in2_valid;
	wire [0 : 0]branchC_17_out1_data;
	wire branchC_17_out1_ready;
	wire branchC_17_out1_valid;
	wire [0 : 0]branchC_17_out2_data;
	wire branchC_17_out2_ready;
	wire branchC_17_out2_valid;

	wire source_0_clk;
	wire source_0_rst;
	wire [2 : 0]source_0_out1_data;
	wire source_0_out1_ready;
	wire source_0_out1_valid;

	wire source_1_clk;
	wire source_1_rst;
	wire [2 : 0]source_1_out1_data;
	wire source_1_out1_ready;
	wire source_1_out1_valid;

	wire source_2_clk;
	wire source_2_rst;
	wire [0 : 0]source_2_out1_data;
	wire source_2_out1_ready;
	wire source_2_out1_valid;

	wire source_3_clk;
	wire source_3_rst;
	wire [5 : 0]source_3_out1_data;
	wire source_3_out1_ready;
	wire source_3_out1_valid;

	wire fork_27_clk;
	wire fork_27_rst;
	wire [0 : 0]fork_27_in1_data;
	wire fork_27_in1_ready;
	wire fork_27_in1_valid;
	wire [0 : 0]fork_27_out1_data;
	wire fork_27_out1_ready;
	wire fork_27_out1_valid;
	wire [0 : 0]fork_27_out2_data;
	wire fork_27_out2_ready;
	wire fork_27_out2_valid;

	wire cst_8_clk;
	wire cst_8_rst;
	wire [2 : 0]cst_8_in1_data;
	wire cst_8_in1_ready;
	wire cst_8_in1_valid;
	wire [2 : 0]cst_8_out1_data;
	wire cst_8_out1_ready;
	wire cst_8_out1_valid;

	wire shl_22_clk;
	wire shl_22_rst;
	wire [10 : 0]shl_22_in1_data;
	wire shl_22_in1_ready;
	wire shl_22_in1_valid;
	wire [10 : 0]shl_22_in2_data;
	wire shl_22_in2_ready;
	wire shl_22_in2_valid;
	wire [10 : 0]shl_22_out1_data;
	wire shl_22_out1_ready;
	wire shl_22_out1_valid;

	wire add_23_clk;
	wire add_23_rst;
	wire [11 : 0]add_23_in1_data;
	wire add_23_in1_ready;
	wire add_23_in1_valid;
	wire [11 : 0]add_23_in2_data;
	wire add_23_in2_ready;
	wire add_23_in2_valid;
	wire [11 : 0]add_23_out1_data;
	wire add_23_out1_ready;
	wire add_23_out1_valid;

	wire store_0_clk;
	wire store_0_rst;
	wire [31 : 0]store_0_in1_data;
	wire store_0_in1_ready;
	wire store_0_in1_valid;
	wire [11 : 0]store_0_in2_data;
	wire store_0_in2_ready;
	wire store_0_in2_valid;
	wire [31 : 0]store_0_out1_data;
	wire store_0_out1_ready;
	wire store_0_out1_valid;
	wire [11 : 0]store_0_out2_data;
	wire store_0_out2_ready;
	wire store_0_out2_valid;

	wire cst_9_clk;
	wire cst_9_rst;
	wire [0 : 0]cst_9_in1_data;
	wire cst_9_in1_ready;
	wire cst_9_in1_valid;
	wire [0 : 0]cst_9_out1_data;
	wire cst_9_out1_ready;
	wire cst_9_out1_valid;

	wire add_26_clk;
	wire add_26_rst;
	wire [5 : 0]add_26_in1_data;
	wire add_26_in1_ready;
	wire add_26_in1_valid;
	wire [5 : 0]add_26_in2_data;
	wire add_26_in2_ready;
	wire add_26_in2_valid;
	wire [5 : 0]add_26_out1_data;
	wire add_26_out1_ready;
	wire add_26_out1_valid;

	wire cst_10_clk;
	wire cst_10_rst;
	wire [5 : 0]cst_10_in1_data;
	wire cst_10_in1_ready;
	wire cst_10_in1_valid;
	wire [5 : 0]cst_10_out1_data;
	wire cst_10_out1_ready;
	wire cst_10_out1_valid;

	wire icmp_27_clk;
	wire icmp_27_rst;
	wire [5 : 0]icmp_27_in1_data;
	wire icmp_27_in1_ready;
	wire icmp_27_in1_valid;
	wire [5 : 0]icmp_27_in2_data;
	wire icmp_27_in2_ready;
	wire icmp_27_in2_valid;
	wire [0 : 0]icmp_27_out1_data;
	wire icmp_27_out1_ready;
	wire icmp_27_out1_valid;

	wire phi_n2_clk;
	wire phi_n2_rst;
	wire [5 : 0]phi_n2_in1_data;
	wire phi_n2_in1_ready;
	wire phi_n2_in1_valid;
	wire [5 : 0]phi_n2_out1_data;
	wire phi_n2_out1_ready;
	wire phi_n2_out1_valid;

	wire phi_n3_clk;
	wire phi_n3_rst;
	wire [5 : 0]phi_n3_in1_data;
	wire phi_n3_in1_ready;
	wire phi_n3_in1_valid;
	wire [5 : 0]phi_n3_out1_data;
	wire phi_n3_out1_ready;
	wire phi_n3_out1_valid;

	wire phi_n4_clk;
	wire phi_n4_rst;
	wire [31 : 0]phi_n4_in1_data;
	wire phi_n4_in1_ready;
	wire phi_n4_in1_valid;
	wire [31 : 0]phi_n4_out1_data;
	wire phi_n4_out1_ready;
	wire phi_n4_out1_valid;

	wire fork_3_clk;
	wire fork_3_rst;
	wire [5 : 0]fork_3_in1_data;
	wire fork_3_in1_ready;
	wire fork_3_in1_valid;
	wire [5 : 0]fork_3_out1_data;
	wire fork_3_out1_ready;
	wire fork_3_out1_valid;
	wire [5 : 0]fork_3_out2_data;
	wire fork_3_out2_ready;
	wire fork_3_out2_valid;

	wire fork_5_clk;
	wire fork_5_rst;
	wire [5 : 0]fork_5_in1_data;
	wire fork_5_in1_ready;
	wire fork_5_in1_valid;
	wire [5 : 0]fork_5_out1_data;
	wire fork_5_out1_ready;
	wire fork_5_out1_valid;
	wire [5 : 0]fork_5_out2_data;
	wire fork_5_out2_ready;
	wire fork_5_out2_valid;

	wire fork_6_clk;
	wire fork_6_rst;
	wire [5 : 0]fork_6_in1_data;
	wire fork_6_in1_ready;
	wire fork_6_in1_valid;
	wire [5 : 0]fork_6_out1_data;
	wire fork_6_out1_ready;
	wire fork_6_out1_valid;
	wire [5 : 0]fork_6_out2_data;
	wire fork_6_out2_ready;
	wire fork_6_out2_valid;

	wire branch_11_clk;
	wire branch_11_rst;
	wire [5 : 0]branch_11_in1_data;
	wire branch_11_in1_ready;
	wire branch_11_in1_valid;
	wire [0 : 0]branch_11_in2_data;
	wire branch_11_in2_ready;
	wire branch_11_in2_valid;
	wire [5 : 0]branch_11_out1_data;
	wire branch_11_out1_ready;
	wire branch_11_out1_valid;
	wire [5 : 0]branch_11_out2_data;
	wire branch_11_out2_ready;
	wire branch_11_out2_valid;

	wire branch_12_clk;
	wire branch_12_rst;
	wire [5 : 0]branch_12_in1_data;
	wire branch_12_in1_ready;
	wire branch_12_in1_valid;
	wire [0 : 0]branch_12_in2_data;
	wire branch_12_in2_ready;
	wire branch_12_in2_valid;
	wire [5 : 0]branch_12_out1_data;
	wire branch_12_out1_ready;
	wire branch_12_out1_valid;
	wire [5 : 0]branch_12_out2_data;
	wire branch_12_out2_ready;
	wire branch_12_out2_valid;

	wire fork_13_clk;
	wire fork_13_rst;
	wire [0 : 0]fork_13_in1_data;
	wire fork_13_in1_ready;
	wire fork_13_in1_valid;
	wire [0 : 0]fork_13_out1_data;
	wire fork_13_out1_ready;
	wire fork_13_out1_valid;
	wire [0 : 0]fork_13_out2_data;
	wire fork_13_out2_ready;
	wire fork_13_out2_valid;
	wire [0 : 0]fork_13_out3_data;
	wire fork_13_out3_ready;
	wire fork_13_out3_valid;

	wire cst_13_clk;
	wire cst_13_rst;
	wire [0 : 0]cst_13_in1_data;
	wire cst_13_in1_ready;
	wire cst_13_in1_valid;
	wire [0 : 0]cst_13_out1_data;
	wire cst_13_out1_ready;
	wire cst_13_out1_valid;

	wire phiC_10_clk;
	wire phiC_10_rst;
	wire [0 : 0]phiC_10_in1_data;
	wire phiC_10_in1_ready;
	wire phiC_10_in1_valid;
	wire [0 : 0]phiC_10_out1_data;
	wire phiC_10_out1_ready;
	wire phiC_10_out1_valid;

	wire forkC_21_clk;
	wire forkC_21_rst;
	wire [0 : 0]forkC_21_in1_data;
	wire forkC_21_in1_ready;
	wire forkC_21_in1_valid;
	wire [0 : 0]forkC_21_out1_data;
	wire forkC_21_out1_ready;
	wire forkC_21_out1_valid;
	wire [0 : 0]forkC_21_out2_data;
	wire forkC_21_out2_ready;
	wire forkC_21_out2_valid;

	wire branchC_18_clk;
	wire branchC_18_rst;
	wire [0 : 0]branchC_18_in1_data;
	wire branchC_18_in1_ready;
	wire branchC_18_in1_valid;
	wire [0 : 0]branchC_18_in2_data;
	wire branchC_18_in2_ready;
	wire branchC_18_in2_valid;
	wire [0 : 0]branchC_18_out1_data;
	wire branchC_18_out1_ready;
	wire branchC_18_out1_valid;
	wire [0 : 0]branchC_18_out2_data;
	wire branchC_18_out2_ready;
	wire branchC_18_out2_valid;

	wire source_4_clk;
	wire source_4_rst;
	wire [2 : 0]source_4_out1_data;
	wire source_4_out1_ready;
	wire source_4_out1_valid;

	wire source_5_clk;
	wire source_5_rst;
	wire [0 : 0]source_5_out1_data;
	wire source_5_out1_ready;
	wire source_5_out1_valid;

	wire source_6_clk;
	wire source_6_rst;
	wire [5 : 0]source_6_out1_data;
	wire source_6_out1_ready;
	wire source_6_out1_valid;

	wire ret_0_clk;
	wire ret_0_rst;
	wire [0 : 0]ret_0_in1_data;
	wire ret_0_in1_ready;
	wire ret_0_in1_valid;
	wire [0 : 0]ret_0_out1_data;
	wire ret_0_out1_ready;
	wire ret_0_out1_valid;

	wire end_0_clk;
	wire end_0_rst;
	wire [0 : 0]end_0_in1_data;
	wire end_0_in1_ready;
	wire end_0_in1_valid;
	wire [0 : 0]end_0_in2_data;
	wire end_0_in2_ready;
	wire end_0_in2_valid;
	wire [0 : 0]end_0_in3_data;
	wire end_0_in3_ready;
	wire end_0_in3_valid;
	wire [0 : 0]end_0_in4_data;
	wire end_0_in4_ready;
	wire end_0_in4_valid;
	wire [0 : 0]end_0_out1_data;
	wire end_0_out1_ready;
	wire end_0_out1_valid;

	wire phiC_12_clk;
	wire phiC_12_rst;
	wire [0 : 0]phiC_12_in1_data;
	wire phiC_12_in1_ready;
	wire phiC_12_in1_valid;
	wire [0 : 0]phiC_12_out1_data;
	wire phiC_12_out1_ready;
	wire phiC_12_out1_valid;

	wire phi_1_clk;
	wire phi_1_rst;
	wire [0 : 0]phi_1_in1_data;
	wire phi_1_in1_ready;
	wire phi_1_in1_valid;
	wire [5 : 0]phi_1_in2_data;
	wire phi_1_in2_ready;
	wire phi_1_in2_valid;
	wire [5 : 0]phi_1_in3_data;
	wire phi_1_in3_ready;
	wire phi_1_in3_valid;
	wire [5 : 0]phi_1_out1_data;
	wire phi_1_out1_ready;
	wire phi_1_out1_valid;

	wire brCst_block2_clk;
	wire brCst_block2_rst;
	wire [0 : 0]brCst_block2_in1_data;
	wire brCst_block2_in1_ready;
	wire brCst_block2_in1_valid;
	wire [0 : 0]brCst_block2_out1_data;
	wire brCst_block2_out1_ready;
	wire brCst_block2_out1_valid;

	wire cst_1_clk;
	wire cst_1_rst;
	wire [0 : 0]cst_1_in1_data;
	wire cst_1_in1_ready;
	wire cst_1_in1_valid;
	wire [0 : 0]cst_1_out1_data;
	wire cst_1_out1_ready;
	wire cst_1_out1_valid;

	wire branch_1_clk;
	wire branch_1_rst;
	wire [0 : 0]branch_1_in1_data;
	wire branch_1_in1_ready;
	wire branch_1_in1_valid;
	wire [0 : 0]branch_1_in2_data;
	wire branch_1_in2_ready;
	wire branch_1_in2_valid;
	wire [0 : 0]branch_1_out1_data;
	wire branch_1_out1_ready;
	wire branch_1_out1_valid;
	wire [0 : 0]branch_1_out2_data;
	wire branch_1_out2_ready;
	wire branch_1_out2_valid;

	wire branch_2_clk;
	wire branch_2_rst;
	wire [5 : 0]branch_2_in1_data;
	wire branch_2_in1_ready;
	wire branch_2_in1_valid;
	wire [0 : 0]branch_2_in2_data;
	wire branch_2_in2_ready;
	wire branch_2_in2_valid;
	wire [5 : 0]branch_2_out1_data;
	wire branch_2_out1_ready;
	wire branch_2_out1_valid;
	wire [5 : 0]branch_2_out2_data;
	wire branch_2_out2_ready;
	wire branch_2_out2_valid;

	wire fork_10_clk;
	wire fork_10_rst;
	wire [0 : 0]fork_10_in1_data;
	wire fork_10_in1_ready;
	wire fork_10_in1_valid;
	wire [0 : 0]fork_10_out1_data;
	wire fork_10_out1_ready;
	wire fork_10_out1_valid;
	wire [0 : 0]fork_10_out2_data;
	wire fork_10_out2_ready;
	wire fork_10_out2_valid;
	wire [0 : 0]fork_10_out3_data;
	wire fork_10_out3_ready;
	wire fork_10_out3_valid;

	wire phiC_7_clk;
	wire phiC_7_rst;
	wire [0 : 0]phiC_7_in1_data;
	wire phiC_7_in1_ready;
	wire phiC_7_in1_valid;
	wire [0 : 0]phiC_7_in2_data;
	wire phiC_7_in2_ready;
	wire phiC_7_in2_valid;
	wire [0 : 0]phiC_7_out1_data;
	wire phiC_7_out1_ready;
	wire phiC_7_out1_valid;
	wire [0 : 0]phiC_7_out2_data;
	wire phiC_7_out2_ready;
	wire phiC_7_out2_valid;

	wire forkC_18_clk;
	wire forkC_18_rst;
	wire [0 : 0]forkC_18_in1_data;
	wire forkC_18_in1_ready;
	wire forkC_18_in1_valid;
	wire [0 : 0]forkC_18_out1_data;
	wire forkC_18_out1_ready;
	wire forkC_18_out1_valid;
	wire [0 : 0]forkC_18_out2_data;
	wire forkC_18_out2_ready;
	wire forkC_18_out2_valid;
	wire [0 : 0]forkC_18_out3_data;
	wire forkC_18_out3_ready;
	wire forkC_18_out3_valid;

	wire branchC_15_clk;
	wire branchC_15_rst;
	wire [0 : 0]branchC_15_in1_data;
	wire branchC_15_in1_ready;
	wire branchC_15_in1_valid;
	wire [0 : 0]branchC_15_in2_data;
	wire branchC_15_in2_ready;
	wire branchC_15_in2_valid;
	wire [0 : 0]branchC_15_out1_data;
	wire branchC_15_out1_ready;
	wire branchC_15_out1_valid;
	wire [0 : 0]branchC_15_out2_data;
	wire branchC_15_out2_ready;
	wire branchC_15_out2_valid;

	wire MC_in_a_clk;
	wire MC_in_a_rst;
	wire [11 : 0]MC_in_a_in1_data;
	wire MC_in_a_in1_ready;
	wire MC_in_a_in1_valid;
	wire [31 : 0]MC_in_a_in2_data;
	wire MC_in_a_in2_ready;
	wire MC_in_a_in2_valid;
	wire [11 : 0]MC_in_a_in3_data;
	wire MC_in_a_in3_ready;
	wire MC_in_a_in3_valid;
	wire [31 : 0]MC_in_a_in4_data;
	wire MC_in_a_in4_ready;
	wire MC_in_a_in4_valid;
	wire [31 : 0]MC_in_a_out1_data;
	wire MC_in_a_out1_ready;
	wire MC_in_a_out1_valid;
	wire [0 : 0]MC_in_a_out2_data;
	wire MC_in_a_out2_ready;
	wire MC_in_a_out2_valid;

	wire MC_in_b_clk;
	wire MC_in_b_rst;
	wire [11 : 0]MC_in_b_in1_data;
	wire MC_in_b_in1_ready;
	wire MC_in_b_in1_valid;
	wire [31 : 0]MC_in_b_in2_data;
	wire MC_in_b_in2_ready;
	wire MC_in_b_in2_valid;
	wire [11 : 0]MC_in_b_in3_data;
	wire MC_in_b_in3_ready;
	wire MC_in_b_in3_valid;
	wire [31 : 0]MC_in_b_in4_data;
	wire MC_in_b_in4_ready;
	wire MC_in_b_in4_valid;
	wire [31 : 0]MC_in_b_out1_data;
	wire MC_in_b_out1_ready;
	wire MC_in_b_out1_valid;
	wire [0 : 0]MC_in_b_out2_data;
	wire MC_in_b_out2_ready;
	wire MC_in_b_out2_valid;

	wire MC_out_c_clk;
	wire MC_out_c_rst;
	wire [31 : 0]MC_out_c_in1_data;
	wire MC_out_c_in1_ready;
	wire MC_out_c_in1_valid;
	wire [11 : 0]MC_out_c_in2_data;
	wire MC_out_c_in2_ready;
	wire MC_out_c_in2_valid;
	wire [31 : 0]MC_out_c_in3_data;
	wire MC_out_c_in3_ready;
	wire MC_out_c_in3_valid;
	wire [11 : 0]MC_out_c_in4_data;
	wire MC_out_c_in4_ready;
	wire MC_out_c_in4_valid;
	wire [0 : 0]MC_out_c_out1_data;
	wire MC_out_c_out1_ready;
	wire MC_out_c_out1_valid;
	wire [31 : 0]MC_out_c_out2_data;
	wire MC_out_c_out2_ready;
	wire MC_out_c_out2_valid;

	wire sink_0_clk;
	wire sink_0_rst;
	wire [0 : 0]sink_0_in1_data;
	wire sink_0_in1_ready;
	wire sink_0_in1_valid;

	wire sink_1_clk;
	wire sink_1_rst;
	wire [0 : 0]sink_1_in1_data;
	wire sink_1_in1_ready;
	wire sink_1_in1_valid;

	wire sink_2_clk;
	wire sink_2_rst;
	wire [5 : 0]sink_2_in1_data;
	wire sink_2_in1_ready;
	wire sink_2_in1_valid;

	wire sink_3_clk;
	wire sink_3_rst;
	wire [0 : 0]sink_3_in1_data;
	wire sink_3_in1_ready;
	wire sink_3_in1_valid;

	wire sink_4_clk;
	wire sink_4_rst;
	wire [0 : 0]sink_4_in1_data;
	wire sink_4_in1_ready;
	wire sink_4_in1_valid;

	wire sink_5_clk;
	wire sink_5_rst;
	wire [5 : 0]sink_5_in1_data;
	wire sink_5_in1_ready;
	wire sink_5_in1_valid;

	wire sink_6_clk;
	wire sink_6_rst;
	wire [5 : 0]sink_6_in1_data;
	wire sink_6_in1_ready;
	wire sink_6_in1_valid;

	wire sink_7_clk;
	wire sink_7_rst;
	wire [5 : 0]sink_7_in1_data;
	wire sink_7_in1_ready;
	wire sink_7_in1_valid;

	wire sink_8_clk;
	wire sink_8_rst;
	wire [5 : 0]sink_8_in1_data;
	wire sink_8_in1_ready;
	wire sink_8_in1_valid;

	wire sink_9_clk;
	wire sink_9_rst;
	wire [5 : 0]sink_9_in1_data;
	wire sink_9_in1_ready;
	wire sink_9_in1_valid;

	wire sink_10_clk;
	wire sink_10_rst;
	wire [0 : 0]sink_10_in1_data;
	wire sink_10_in1_ready;
	wire sink_10_in1_valid;

	wire sink_11_clk;
	wire sink_11_rst;
	wire [0 : 0]sink_11_in1_data;
	wire sink_11_in1_ready;
	wire sink_11_in1_valid;

	wire sink_12_clk;
	wire sink_12_rst;
	wire [0 : 0]sink_12_in1_data;
	wire sink_12_in1_ready;
	wire sink_12_in1_valid;

	wire Buffer_100_clk;
	wire Buffer_100_rst;
	wire [31 : 0]Buffer_100_in1_data;
	wire Buffer_100_in1_ready;
	wire Buffer_100_in1_valid;
	wire [31 : 0]Buffer_100_out1_data;
	wire Buffer_100_out1_ready;
	wire Buffer_100_out1_valid;

	wire Buffer_101_clk;
	wire Buffer_101_rst;
	wire [31 : 0]Buffer_101_in1_data;
	wire Buffer_101_in1_ready;
	wire Buffer_101_in1_valid;
	wire [31 : 0]Buffer_101_out1_data;
	wire Buffer_101_out1_ready;
	wire Buffer_101_out1_valid;

	wire Buffer_102_clk;
	wire Buffer_102_rst;
	wire [31 : 0]Buffer_102_in1_data;
	wire Buffer_102_in1_ready;
	wire Buffer_102_in1_valid;
	wire [31 : 0]Buffer_102_out1_data;
	wire Buffer_102_out1_ready;
	wire Buffer_102_out1_valid;

	wire Buffer_103_clk;
	wire Buffer_103_rst;
	wire [31 : 0]Buffer_103_in1_data;
	wire Buffer_103_in1_ready;
	wire Buffer_103_in1_valid;
	wire [31 : 0]Buffer_103_out1_data;
	wire Buffer_103_out1_ready;
	wire Buffer_103_out1_valid;

	wire Buffer_104_clk;
	wire Buffer_104_rst;
	wire [31 : 0]Buffer_104_in1_data;
	wire Buffer_104_in1_ready;
	wire Buffer_104_in1_valid;
	wire [31 : 0]Buffer_104_out1_data;
	wire Buffer_104_out1_ready;
	wire Buffer_104_out1_valid;

	wire Buffer_105_clk;
	wire Buffer_105_rst;
	wire [31 : 0]Buffer_105_in1_data;
	wire Buffer_105_in1_ready;
	wire Buffer_105_in1_valid;
	wire [31 : 0]Buffer_105_out1_data;
	wire Buffer_105_out1_ready;
	wire Buffer_105_out1_valid;

	wire Buffer_106_clk;
	wire Buffer_106_rst;
	wire [31 : 0]Buffer_106_in1_data;
	wire Buffer_106_in1_ready;
	wire Buffer_106_in1_valid;
	wire [31 : 0]Buffer_106_out1_data;
	wire Buffer_106_out1_ready;
	wire Buffer_106_out1_valid;

	wire Buffer_107_clk;
	wire Buffer_107_rst;
	wire [31 : 0]Buffer_107_in1_data;
	wire Buffer_107_in1_ready;
	wire Buffer_107_in1_valid;
	wire [31 : 0]Buffer_107_out1_data;
	wire Buffer_107_out1_ready;
	wire Buffer_107_out1_valid;

	wire Buffer_108_clk;
	wire Buffer_108_rst;
	wire [31 : 0]Buffer_108_in1_data;
	wire Buffer_108_in1_ready;
	wire Buffer_108_in1_valid;
	wire [31 : 0]Buffer_108_out1_data;
	wire Buffer_108_out1_ready;
	wire Buffer_108_out1_valid;

	wire Buffer_109_clk;
	wire Buffer_109_rst;
	wire [31 : 0]Buffer_109_in1_data;
	wire Buffer_109_in1_ready;
	wire Buffer_109_in1_valid;
	wire [31 : 0]Buffer_109_out1_data;
	wire Buffer_109_out1_ready;
	wire Buffer_109_out1_valid;



	assign brCst_block1_clk = clk;
	assign brCst_block1_rst = rst;
	assign fork_17_in1_data = brCst_block1_out1_data;
	assign fork_17_in1_valid = brCst_block1_out1_valid;
	assign brCst_block1_out1_ready = fork_17_in1_ready;

	assign cst_0_clk = clk;
	assign cst_0_rst = rst;
	assign branch_0_in1_data = cst_0_out1_data;
	assign branch_0_in1_valid = cst_0_out1_valid;
	assign cst_0_out1_ready = branch_0_in1_ready;

	assign branch_0_clk = clk;
	assign branch_0_rst = rst;
	assign phi_1_in2_data = branch_0_out1_data;
	assign phi_1_in2_valid = branch_0_out1_valid;
	assign branch_0_out1_ready = phi_1_in2_ready;
	assign sink_0_in1_data = branch_0_out2_data;
	assign sink_0_in1_valid = branch_0_out2_valid;
	assign branch_0_out2_ready = sink_0_in1_ready;

	assign start_0_clk = clk;
	assign start_0_rst = rst;
	assign start_0_in1_data = start_in;
	assign start_0_in1_valid = start_valid;
	assign start_ready = start_0_in1_ready;
	assign forkC_16_in1_data = start_0_out1_data;
	assign forkC_16_in1_valid = start_0_out1_valid;
	assign start_0_out1_ready = forkC_16_in1_ready;

	assign forkC_16_clk = clk;
	assign forkC_16_rst = rst;
	assign cst_0_in1_data = forkC_16_out1_data;
	assign cst_0_in1_valid = forkC_16_out1_valid;
	assign forkC_16_out1_ready = cst_0_in1_ready;
	assign branchC_14_in1_data = forkC_16_out2_data;
	assign branchC_14_in1_valid = forkC_16_out2_valid;
	assign forkC_16_out2_ready = branchC_14_in1_ready;
	assign brCst_block1_in1_data = forkC_16_out3_data;
	assign brCst_block1_in1_valid = forkC_16_out3_valid;
	assign forkC_16_out3_ready = brCst_block1_in1_ready;

	assign branchC_14_clk = clk;
	assign branchC_14_rst = rst;
	assign phiC_7_in1_data = branchC_14_out1_data;
	assign phiC_7_in1_valid = branchC_14_out1_valid;
	assign branchC_14_out1_ready = phiC_7_in1_ready;
	assign sink_10_in1_data = branchC_14_out2_data;
	assign sink_10_in1_valid = branchC_14_out2_valid;
	assign branchC_14_out2_ready = sink_10_in1_ready;

	assign fork_17_clk = clk;
	assign fork_17_rst = rst;
	assign branch_0_in2_data = fork_17_out1_data;
	assign branch_0_in2_valid = fork_17_out1_valid;
	assign fork_17_out1_ready = branch_0_in2_ready;
	assign branchC_14_in2_data = fork_17_out2_data;
	assign branchC_14_in2_valid = fork_17_out2_valid;
	assign fork_17_out2_ready = branchC_14_in2_ready;

	assign phi_3_clk = clk;
	assign phi_3_rst = rst;
	assign branch_5_in1_data = phi_3_out1_data;
	assign branch_5_in1_valid = phi_3_out1_valid;
	assign phi_3_out1_ready = branch_5_in1_ready;

	assign brCst_block3_clk = clk;
	assign brCst_block3_rst = rst;
	assign fork_11_in1_data = brCst_block3_out1_data;
	assign fork_11_in1_valid = brCst_block3_out1_valid;
	assign brCst_block3_out1_ready = fork_11_in1_ready;

	assign cst_2_clk = clk;
	assign cst_2_rst = rst;
	assign branch_3_in1_data = cst_2_out1_data;
	assign branch_3_in1_valid = cst_2_out1_valid;
	assign cst_2_out1_ready = branch_3_in1_ready;

	assign cst_3_clk = clk;
	assign cst_3_rst = rst;
	assign branch_4_in1_data = cst_3_out1_data;
	assign branch_4_in1_valid = cst_3_out1_valid;
	assign cst_3_out1_ready = branch_4_in1_ready;

	assign phi_n1_clk = clk;
	assign phi_n1_rst = rst;
	assign branch_6_in1_data = phi_n1_out1_data;
	assign branch_6_in1_valid = phi_n1_out1_valid;
	assign phi_n1_out1_ready = branch_6_in1_ready;

	assign branch_3_clk = clk;
	assign branch_3_rst = rst;
	assign phi_5_in2_data = branch_3_out1_data;
	assign phi_5_in2_valid = branch_3_out1_valid;
	assign branch_3_out1_ready = phi_5_in2_ready;
	assign sink_3_in1_data = branch_3_out2_data;
	assign sink_3_in1_valid = branch_3_out2_valid;
	assign branch_3_out2_ready = sink_3_in1_ready;

	assign branch_4_clk = clk;
	assign branch_4_rst = rst;
	assign phi_6_in2_data = branch_4_out1_data;
	assign phi_6_in2_valid = branch_4_out1_valid;
	assign branch_4_out1_ready = phi_6_in2_ready;
	assign sink_4_in1_data = branch_4_out2_data;
	assign sink_4_in1_valid = branch_4_out2_valid;
	assign branch_4_out2_ready = sink_4_in1_ready;

	assign branch_5_clk = clk;
	assign branch_5_rst = rst;
	assign phi_n6_in1_data = branch_5_out1_data;
	assign phi_n6_in1_valid = branch_5_out1_valid;
	assign branch_5_out1_ready = phi_n6_in1_ready;
	assign sink_5_in1_data = branch_5_out2_data;
	assign sink_5_in1_valid = branch_5_out2_valid;
	assign branch_5_out2_ready = sink_5_in1_ready;

	assign branch_6_clk = clk;
	assign branch_6_rst = rst;
	assign phi_n5_in1_data = branch_6_out1_data;
	assign phi_n5_in1_valid = branch_6_out1_valid;
	assign branch_6_out1_ready = phi_n5_in1_ready;
	assign sink_6_in1_data = branch_6_out2_data;
	assign sink_6_in1_valid = branch_6_out2_valid;
	assign branch_6_out2_ready = sink_6_in1_ready;

	assign fork_11_clk = clk;
	assign fork_11_rst = rst;
	assign branch_6_in2_data = fork_11_out1_data;
	assign branch_6_in2_valid = fork_11_out1_valid;
	assign fork_11_out1_ready = branch_6_in2_ready;
	assign branch_5_in2_data = fork_11_out2_data;
	assign branch_5_in2_valid = fork_11_out2_valid;
	assign fork_11_out2_ready = branch_5_in2_ready;
	assign branch_4_in2_data = fork_11_out3_data;
	assign branch_4_in2_valid = fork_11_out3_valid;
	assign fork_11_out3_ready = branch_4_in2_ready;
	assign branch_3_in2_data = fork_11_out4_data;
	assign branch_3_in2_valid = fork_11_out4_valid;
	assign fork_11_out4_ready = branch_3_in2_ready;
	assign branchC_16_in2_data = fork_11_out5_data;
	assign branchC_16_in2_valid = fork_11_out5_valid;
	assign fork_11_out5_ready = branchC_16_in2_ready;

	assign phiC_8_clk = clk;
	assign phiC_8_rst = rst;
	assign forkC_19_in1_data = phiC_8_out1_data;
	assign forkC_19_in1_valid = phiC_8_out1_valid;
	assign phiC_8_out1_ready = forkC_19_in1_ready;
	assign phi_3_in1_data = phiC_8_out2_data;
	assign phi_3_in1_valid = phiC_8_out2_valid;
	assign phiC_8_out2_ready = phi_3_in1_ready;

	assign forkC_19_clk = clk;
	assign forkC_19_rst = rst;
	assign cst_2_in1_data = forkC_19_out1_data;
	assign cst_2_in1_valid = forkC_19_out1_valid;
	assign forkC_19_out1_ready = cst_2_in1_ready;
	assign cst_3_in1_data = forkC_19_out2_data;
	assign cst_3_in1_valid = forkC_19_out2_valid;
	assign forkC_19_out2_ready = cst_3_in1_ready;
	assign branchC_16_in1_data = forkC_19_out3_data;
	assign branchC_16_in1_valid = forkC_19_out3_valid;
	assign forkC_19_out3_ready = branchC_16_in1_ready;
	assign brCst_block3_in1_data = forkC_19_out4_data;
	assign brCst_block3_in1_valid = forkC_19_out4_valid;
	assign forkC_19_out4_ready = brCst_block3_in1_ready;

	assign branchC_16_clk = clk;
	assign branchC_16_rst = rst;
	assign phiC_9_in1_data = branchC_16_out1_data;
	assign phiC_9_in1_valid = branchC_16_out1_valid;
	assign branchC_16_out1_ready = phiC_9_in1_ready;
	assign sink_12_in1_data = branchC_16_out2_data;
	assign sink_12_in1_valid = branchC_16_out2_valid;
	assign branchC_16_out2_ready = sink_12_in1_ready;

	assign cst_11_clk = clk;
	assign cst_11_rst = rst;
	assign add_29_in2_data = cst_11_out1_data;
	assign add_29_in2_valid = cst_11_out1_valid;
	assign cst_11_out1_ready = add_29_in2_ready;

	assign add_29_clk = clk;
	assign add_29_rst = rst;
	assign fork_4_in1_data = add_29_out1_data;
	assign fork_4_in1_valid = add_29_out1_valid;
	assign add_29_out1_ready = fork_4_in1_ready;

	assign cst_12_clk = clk;
	assign cst_12_rst = rst;
	assign icmp_30_in2_data = cst_12_out1_data;
	assign icmp_30_in2_valid = cst_12_out1_valid;
	assign cst_12_out1_ready = icmp_30_in2_ready;

	assign icmp_30_clk = clk;
	assign icmp_30_rst = rst;
	assign fork_23_in1_data = icmp_30_out1_data;
	assign fork_23_in1_valid = icmp_30_out1_valid;
	assign icmp_30_out1_ready = fork_23_in1_ready;

	assign phi_n0_clk = clk;
	assign phi_n0_rst = rst;
	assign add_29_in1_data = phi_n0_out1_data;
	assign add_29_in1_valid = phi_n0_out1_valid;
	assign phi_n0_out1_ready = add_29_in1_ready;

	assign fork_4_clk = clk;
	assign fork_4_rst = rst;
	assign icmp_30_in1_data = fork_4_out1_data;
	assign icmp_30_in1_valid = fork_4_out1_valid;
	assign fork_4_out1_ready = icmp_30_in1_ready;
	assign branch_13_in1_data = fork_4_out2_data;
	assign branch_13_in1_valid = fork_4_out2_valid;
	assign fork_4_out2_ready = branch_13_in1_ready;

	assign branch_13_clk = clk;
	assign branch_13_rst = rst;
	assign Buffer_108_in1_data = branch_13_out1_data;
	assign Buffer_108_in1_valid = branch_13_out1_valid;
	assign branch_13_out1_ready = Buffer_108_in1_ready;
	assign sink_9_in1_data = branch_13_out2_data;
	assign sink_9_in1_valid = branch_13_out2_valid;
	assign branch_13_out2_ready = sink_9_in1_ready;

	assign phiC_11_clk = clk;
	assign phiC_11_rst = rst;
	assign branchC_19_in1_data = phiC_11_out1_data;
	assign branchC_19_in1_valid = phiC_11_out1_valid;
	assign phiC_11_out1_ready = branchC_19_in1_ready;

	assign branchC_19_clk = clk;
	assign branchC_19_rst = rst;
	assign Buffer_109_in1_data = branchC_19_out1_data;
	assign Buffer_109_in1_valid = branchC_19_out1_valid;
	assign branchC_19_out1_ready = Buffer_109_in1_ready;
	assign phiC_12_in1_data = branchC_19_out2_data;
	assign phiC_12_in1_valid = branchC_19_out2_valid;
	assign branchC_19_out2_ready = phiC_12_in1_ready;

	assign fork_23_clk = clk;
	assign fork_23_rst = rst;
	assign branch_13_in2_data = fork_23_out1_data;
	assign branch_13_in2_valid = fork_23_out1_valid;
	assign fork_23_out1_ready = branch_13_in2_ready;
	assign branchC_19_in2_data = fork_23_out2_data;
	assign branchC_19_in2_valid = fork_23_out2_valid;
	assign fork_23_out2_ready = branchC_19_in2_ready;

	assign source_7_clk = clk;
	assign source_7_rst = rst;
	assign cst_11_in1_data = source_7_out1_data;
	assign cst_11_in1_valid = source_7_out1_valid;
	assign source_7_out1_ready = cst_11_in1_ready;

	assign source_8_clk = clk;
	assign source_8_rst = rst;
	assign cst_12_in1_data = source_8_out1_data;
	assign cst_12_in1_valid = source_8_out1_valid;
	assign source_8_out1_ready = cst_12_in1_ready;

	assign phi_5_clk = clk;
	assign phi_5_rst = rst;
	assign add_18_in1_data = phi_5_out1_data;
	assign add_18_in1_valid = phi_5_out1_valid;
	assign phi_5_out1_ready = add_18_in1_ready;

	assign phi_6_clk = clk;
	assign phi_6_rst = rst;
	assign fork_0_in1_data = phi_6_out1_data;
	assign fork_0_in1_valid = phi_6_out1_valid;
	assign phi_6_out1_ready = fork_0_in1_ready;

	assign cst_4_clk = clk;
	assign cst_4_rst = rst;
	assign shl_7_in2_data = cst_4_out1_data;
	assign shl_7_in2_valid = cst_4_out1_valid;
	assign cst_4_out1_ready = shl_7_in2_ready;

	assign shl_7_clk = clk;
	assign shl_7_rst = rst;
	assign add_8_in1_data = shl_7_out1_data;
	assign add_8_in1_valid = shl_7_out1_valid;
	assign shl_7_out1_ready = add_8_in1_ready;

	assign add_8_clk = clk;
	assign add_8_rst = rst;
	assign load_11_in2_data = add_8_out1_data;
	assign load_11_in2_valid = add_8_out1_valid;
	assign add_8_out1_ready = load_11_in2_ready;

	assign load_11_clk = clk;
	assign load_11_rst = rst;
	assign mul_17_in1_data = load_11_out1_data;
	assign mul_17_in1_valid = load_11_out1_valid;
	assign load_11_out1_ready = mul_17_in1_ready;
	assign MC_in_a_in1_data = load_11_out2_data;
	assign MC_in_a_in1_valid = load_11_out2_valid;
	assign load_11_out2_ready = MC_in_a_in1_ready;

	assign cst_5_clk = clk;
	assign cst_5_rst = rst;
	assign shl_12_in2_data = cst_5_out1_data;
	assign shl_12_in2_valid = cst_5_out1_valid;
	assign cst_5_out1_ready = shl_12_in2_ready;

	assign shl_12_clk = clk;
	assign shl_12_rst = rst;
	assign add_13_in1_data = shl_12_out1_data;
	assign add_13_in1_valid = shl_12_out1_valid;
	assign shl_12_out1_ready = add_13_in1_ready;

	assign add_13_clk = clk;
	assign add_13_rst = rst;
	assign load_16_in2_data = add_13_out1_data;
	assign load_16_in2_valid = add_13_out1_valid;
	assign add_13_out1_ready = load_16_in2_ready;

	assign load_16_clk = clk;
	assign load_16_rst = rst;
	assign mul_17_in2_data = load_16_out1_data;
	assign mul_17_in2_valid = load_16_out1_valid;
	assign load_16_out1_ready = mul_17_in2_ready;
	assign MC_in_b_in1_data = load_16_out2_data;
	assign MC_in_b_in1_valid = load_16_out2_valid;
	assign load_16_out2_ready = MC_in_b_in1_ready;

	assign mul_17_clk = clk;
	assign mul_17_rst = rst;
	assign add_18_in2_data = mul_17_out1_data;
	assign add_18_in2_valid = mul_17_out1_valid;
	assign mul_17_out1_ready = add_18_in2_ready;

	assign add_18_clk = clk;
	assign add_18_rst = rst;
	assign branch_7_in1_data = add_18_out1_data;
	assign branch_7_in1_valid = add_18_out1_valid;
	assign add_18_out1_ready = branch_7_in1_ready;

	assign cst_6_clk = clk;
	assign cst_6_rst = rst;
	assign add_19_in2_data = cst_6_out1_data;
	assign add_19_in2_valid = cst_6_out1_valid;
	assign cst_6_out1_ready = add_19_in2_ready;

	assign add_19_clk = clk;
	assign add_19_rst = rst;
	assign fork_2_in1_data = add_19_out1_data;
	assign fork_2_in1_valid = add_19_out1_valid;
	assign add_19_out1_ready = fork_2_in1_ready;

	assign cst_7_clk = clk;
	assign cst_7_rst = rst;
	assign icmp_20_in2_data = cst_7_out1_data;
	assign icmp_20_in2_valid = cst_7_out1_valid;
	assign cst_7_out1_ready = icmp_20_in2_ready;

	assign icmp_20_clk = clk;
	assign icmp_20_rst = rst;
	assign fork_12_in1_data = icmp_20_out1_data;
	assign fork_12_in1_valid = icmp_20_out1_valid;
	assign icmp_20_out1_ready = fork_12_in1_ready;

	assign phi_n5_clk = clk;
	assign phi_n5_rst = rst;
	assign fork_7_in1_data = phi_n5_out1_data;
	assign fork_7_in1_valid = phi_n5_out1_valid;
	assign phi_n5_out1_ready = fork_7_in1_ready;

	assign phi_n6_clk = clk;
	assign phi_n6_rst = rst;
	assign fork_8_in1_data = phi_n6_out1_data;
	assign fork_8_in1_valid = phi_n6_out1_valid;
	assign phi_n6_out1_ready = fork_8_in1_ready;

	assign fork_0_clk = clk;
	assign fork_0_rst = rst;
	assign add_8_in2_data = fork_0_out1_data;
	assign add_8_in2_valid = fork_0_out1_valid;
	assign fork_0_out1_ready = add_8_in2_ready;
	assign shl_12_in1_data = fork_0_out2_data;
	assign shl_12_in1_valid = fork_0_out2_valid;
	assign fork_0_out2_ready = shl_12_in1_ready;
	assign add_19_in1_data = fork_0_out3_data;
	assign add_19_in1_valid = fork_0_out3_valid;
	assign fork_0_out3_ready = add_19_in1_ready;

	assign fork_2_clk = clk;
	assign fork_2_rst = rst;
	assign icmp_20_in1_data = fork_2_out1_data;
	assign icmp_20_in1_valid = fork_2_out1_valid;
	assign fork_2_out1_ready = icmp_20_in1_ready;
	assign branch_8_in1_data = fork_2_out2_data;
	assign branch_8_in1_valid = fork_2_out2_valid;
	assign fork_2_out2_ready = branch_8_in1_ready;

	assign fork_7_clk = clk;
	assign fork_7_rst = rst;
	assign shl_7_in1_data = fork_7_out1_data;
	assign shl_7_in1_valid = fork_7_out1_valid;
	assign fork_7_out1_ready = shl_7_in1_ready;
	assign branch_9_in1_data = fork_7_out2_data;
	assign branch_9_in1_valid = fork_7_out2_valid;
	assign fork_7_out2_ready = branch_9_in1_ready;

	assign fork_8_clk = clk;
	assign fork_8_rst = rst;
	assign add_13_in2_data = fork_8_out1_data;
	assign add_13_in2_valid = fork_8_out1_valid;
	assign fork_8_out1_ready = add_13_in2_ready;
	assign branch_10_in1_data = fork_8_out2_data;
	assign branch_10_in1_valid = fork_8_out2_valid;
	assign fork_8_out2_ready = branch_10_in1_ready;

	assign branch_7_clk = clk;
	assign branch_7_rst = rst;
	assign Buffer_100_in1_data = branch_7_out1_data;
	assign Buffer_100_in1_valid = branch_7_out1_valid;
	assign branch_7_out1_ready = Buffer_100_in1_ready;
	assign phi_n4_in1_data = branch_7_out2_data;
	assign phi_n4_in1_valid = branch_7_out2_valid;
	assign branch_7_out2_ready = phi_n4_in1_ready;

	assign branch_8_clk = clk;
	assign branch_8_rst = rst;
	assign Buffer_101_in1_data = branch_8_out1_data;
	assign Buffer_101_in1_valid = branch_8_out1_valid;
	assign branch_8_out1_ready = Buffer_101_in1_ready;
	assign sink_7_in1_data = branch_8_out2_data;
	assign sink_7_in1_valid = branch_8_out2_valid;
	assign branch_8_out2_ready = sink_7_in1_ready;

	assign branch_9_clk = clk;
	assign branch_9_rst = rst;
	assign Buffer_102_in1_data = branch_9_out1_data;
	assign Buffer_102_in1_valid = branch_9_out1_valid;
	assign branch_9_out1_ready = Buffer_102_in1_ready;
	assign phi_n2_in1_data = branch_9_out2_data;
	assign phi_n2_in1_valid = branch_9_out2_valid;
	assign branch_9_out2_ready = phi_n2_in1_ready;

	assign branch_10_clk = clk;
	assign branch_10_rst = rst;
	assign Buffer_103_in1_data = branch_10_out1_data;
	assign Buffer_103_in1_valid = branch_10_out1_valid;
	assign branch_10_out1_ready = Buffer_103_in1_ready;
	assign phi_n3_in1_data = branch_10_out2_data;
	assign phi_n3_in1_valid = branch_10_out2_valid;
	assign branch_10_out2_ready = phi_n3_in1_ready;

	assign fork_12_clk = clk;
	assign fork_12_rst = rst;
	assign branch_10_in2_data = fork_12_out1_data;
	assign branch_10_in2_valid = fork_12_out1_valid;
	assign fork_12_out1_ready = branch_10_in2_ready;
	assign branch_9_in2_data = fork_12_out2_data;
	assign branch_9_in2_valid = fork_12_out2_valid;
	assign fork_12_out2_ready = branch_9_in2_ready;
	assign branch_8_in2_data = fork_12_out3_data;
	assign branch_8_in2_valid = fork_12_out3_valid;
	assign fork_12_out3_ready = branch_8_in2_ready;
	assign branch_7_in2_data = fork_12_out4_data;
	assign branch_7_in2_valid = fork_12_out4_valid;
	assign fork_12_out4_ready = branch_7_in2_ready;
	assign branchC_17_in2_data = fork_12_out5_data;
	assign branchC_17_in2_valid = fork_12_out5_valid;
	assign fork_12_out5_ready = branchC_17_in2_ready;

	assign phiC_9_clk = clk;
	assign phiC_9_rst = rst;
	assign branchC_17_in1_data = phiC_9_out1_data;
	assign branchC_17_in1_valid = phiC_9_out1_valid;
	assign phiC_9_out1_ready = branchC_17_in1_ready;
	assign fork_27_in1_data = phiC_9_out2_data;
	assign fork_27_in1_valid = phiC_9_out2_valid;
	assign phiC_9_out2_ready = fork_27_in1_ready;

	assign branchC_17_clk = clk;
	assign branchC_17_rst = rst;
	assign Buffer_104_in1_data = branchC_17_out1_data;
	assign Buffer_104_in1_valid = branchC_17_out1_valid;
	assign branchC_17_out1_ready = Buffer_104_in1_ready;
	assign phiC_10_in1_data = branchC_17_out2_data;
	assign phiC_10_in1_valid = branchC_17_out2_valid;
	assign branchC_17_out2_ready = phiC_10_in1_ready;

	assign source_0_clk = clk;
	assign source_0_rst = rst;
	assign cst_4_in1_data = source_0_out1_data;
	assign cst_4_in1_valid = source_0_out1_valid;
	assign source_0_out1_ready = cst_4_in1_ready;

	assign source_1_clk = clk;
	assign source_1_rst = rst;
	assign cst_5_in1_data = source_1_out1_data;
	assign cst_5_in1_valid = source_1_out1_valid;
	assign source_1_out1_ready = cst_5_in1_ready;

	assign source_2_clk = clk;
	assign source_2_rst = rst;
	assign cst_6_in1_data = source_2_out1_data;
	assign cst_6_in1_valid = source_2_out1_valid;
	assign source_2_out1_ready = cst_6_in1_ready;

	assign source_3_clk = clk;
	assign source_3_rst = rst;
	assign cst_7_in1_data = source_3_out1_data;
	assign cst_7_in1_valid = source_3_out1_valid;
	assign source_3_out1_ready = cst_7_in1_ready;

	assign fork_27_clk = clk;
	assign fork_27_rst = rst;
	assign phi_5_in1_data = fork_27_out1_data;
	assign phi_5_in1_valid = fork_27_out1_valid;
	assign fork_27_out1_ready = phi_5_in1_ready;
	assign phi_6_in1_data = fork_27_out2_data;
	assign phi_6_in1_valid = fork_27_out2_valid;
	assign fork_27_out2_ready = phi_6_in1_ready;

	assign cst_8_clk = clk;
	assign cst_8_rst = rst;
	assign shl_22_in2_data = cst_8_out1_data;
	assign shl_22_in2_valid = cst_8_out1_valid;
	assign cst_8_out1_ready = shl_22_in2_ready;

	assign shl_22_clk = clk;
	assign shl_22_rst = rst;
	assign add_23_in1_data = shl_22_out1_data;
	assign add_23_in1_valid = shl_22_out1_valid;
	assign shl_22_out1_ready = add_23_in1_ready;

	assign add_23_clk = clk;
	assign add_23_rst = rst;
	assign store_0_in2_data = add_23_out1_data;
	assign store_0_in2_valid = add_23_out1_valid;
	assign add_23_out1_ready = store_0_in2_ready;

	assign store_0_clk = clk;
	assign store_0_rst = rst;
	assign MC_out_c_in3_data = store_0_out1_data;
	assign MC_out_c_in3_valid = store_0_out1_valid;
	assign store_0_out1_ready = MC_out_c_in3_ready;
	assign MC_out_c_in2_data = store_0_out2_data;
	assign MC_out_c_in2_valid = store_0_out2_valid;
	assign store_0_out2_ready = MC_out_c_in2_ready;

	assign cst_9_clk = clk;
	assign cst_9_rst = rst;
	assign add_26_in2_data = cst_9_out1_data;
	assign add_26_in2_valid = cst_9_out1_valid;
	assign cst_9_out1_ready = add_26_in2_ready;

	assign add_26_clk = clk;
	assign add_26_rst = rst;
	assign fork_3_in1_data = add_26_out1_data;
	assign fork_3_in1_valid = add_26_out1_valid;
	assign add_26_out1_ready = fork_3_in1_ready;

	assign cst_10_clk = clk;
	assign cst_10_rst = rst;
	assign icmp_27_in2_data = cst_10_out1_data;
	assign icmp_27_in2_valid = cst_10_out1_valid;
	assign cst_10_out1_ready = icmp_27_in2_ready;

	assign icmp_27_clk = clk;
	assign icmp_27_rst = rst;
	assign fork_13_in1_data = icmp_27_out1_data;
	assign fork_13_in1_valid = icmp_27_out1_valid;
	assign icmp_27_out1_ready = fork_13_in1_ready;

	assign phi_n2_clk = clk;
	assign phi_n2_rst = rst;
	assign fork_5_in1_data = phi_n2_out1_data;
	assign fork_5_in1_valid = phi_n2_out1_valid;
	assign phi_n2_out1_ready = fork_5_in1_ready;

	assign phi_n3_clk = clk;
	assign phi_n3_rst = rst;
	assign fork_6_in1_data = phi_n3_out1_data;
	assign fork_6_in1_valid = phi_n3_out1_valid;
	assign phi_n3_out1_ready = fork_6_in1_ready;

	assign phi_n4_clk = clk;
	assign phi_n4_rst = rst;
	assign store_0_in1_data = phi_n4_out1_data;
	assign store_0_in1_valid = phi_n4_out1_valid;
	assign phi_n4_out1_ready = store_0_in1_ready;

	assign fork_3_clk = clk;
	assign fork_3_rst = rst;
	assign icmp_27_in1_data = fork_3_out1_data;
	assign icmp_27_in1_valid = fork_3_out1_valid;
	assign fork_3_out1_ready = icmp_27_in1_ready;
	assign branch_11_in1_data = fork_3_out2_data;
	assign branch_11_in1_valid = fork_3_out2_valid;
	assign fork_3_out2_ready = branch_11_in1_ready;

	assign fork_5_clk = clk;
	assign fork_5_rst = rst;
	assign shl_22_in1_data = fork_5_out1_data;
	assign shl_22_in1_valid = fork_5_out1_valid;
	assign fork_5_out1_ready = shl_22_in1_ready;
	assign branch_12_in1_data = fork_5_out2_data;
	assign branch_12_in1_valid = fork_5_out2_valid;
	assign fork_5_out2_ready = branch_12_in1_ready;

	assign fork_6_clk = clk;
	assign fork_6_rst = rst;
	assign add_23_in2_data = fork_6_out1_data;
	assign add_23_in2_valid = fork_6_out1_valid;
	assign fork_6_out1_ready = add_23_in2_ready;
	assign add_26_in1_data = fork_6_out2_data;
	assign add_26_in1_valid = fork_6_out2_valid;
	assign fork_6_out2_ready = add_26_in1_ready;

	assign branch_11_clk = clk;
	assign branch_11_rst = rst;
	assign Buffer_105_in1_data = branch_11_out1_data;
	assign Buffer_105_in1_valid = branch_11_out1_valid;
	assign branch_11_out1_ready = Buffer_105_in1_ready;
	assign sink_8_in1_data = branch_11_out2_data;
	assign sink_8_in1_valid = branch_11_out2_valid;
	assign branch_11_out2_ready = sink_8_in1_ready;

	assign branch_12_clk = clk;
	assign branch_12_rst = rst;
	assign Buffer_106_in1_data = branch_12_out1_data;
	assign Buffer_106_in1_valid = branch_12_out1_valid;
	assign branch_12_out1_ready = Buffer_106_in1_ready;
	assign phi_n0_in1_data = branch_12_out2_data;
	assign phi_n0_in1_valid = branch_12_out2_valid;
	assign branch_12_out2_ready = phi_n0_in1_ready;

	assign fork_13_clk = clk;
	assign fork_13_rst = rst;
	assign branch_12_in2_data = fork_13_out1_data;
	assign branch_12_in2_valid = fork_13_out1_valid;
	assign fork_13_out1_ready = branch_12_in2_ready;
	assign branch_11_in2_data = fork_13_out2_data;
	assign branch_11_in2_valid = fork_13_out2_valid;
	assign fork_13_out2_ready = branch_11_in2_ready;
	assign branchC_18_in2_data = fork_13_out3_data;
	assign branchC_18_in2_valid = fork_13_out3_valid;
	assign fork_13_out3_ready = branchC_18_in2_ready;

	assign cst_13_clk = clk;
	assign cst_13_rst = rst;
	assign MC_out_c_in1_data = cst_13_out1_data;
	assign MC_out_c_in1_valid = cst_13_out1_valid;
	assign cst_13_out1_ready = MC_out_c_in1_ready;

	assign phiC_10_clk = clk;
	assign phiC_10_rst = rst;
	assign forkC_21_in1_data = phiC_10_out1_data;
	assign forkC_21_in1_valid = phiC_10_out1_valid;
	assign phiC_10_out1_ready = forkC_21_in1_ready;

	assign forkC_21_clk = clk;
	assign forkC_21_rst = rst;
	assign cst_13_in1_data = forkC_21_out1_data;
	assign cst_13_in1_valid = forkC_21_out1_valid;
	assign forkC_21_out1_ready = cst_13_in1_ready;
	assign branchC_18_in1_data = forkC_21_out2_data;
	assign branchC_18_in1_valid = forkC_21_out2_valid;
	assign forkC_21_out2_ready = branchC_18_in1_ready;

	assign branchC_18_clk = clk;
	assign branchC_18_rst = rst;
	assign Buffer_107_in1_data = branchC_18_out1_data;
	assign Buffer_107_in1_valid = branchC_18_out1_valid;
	assign branchC_18_out1_ready = Buffer_107_in1_ready;
	assign phiC_11_in1_data = branchC_18_out2_data;
	assign phiC_11_in1_valid = branchC_18_out2_valid;
	assign branchC_18_out2_ready = phiC_11_in1_ready;

	assign source_4_clk = clk;
	assign source_4_rst = rst;
	assign cst_8_in1_data = source_4_out1_data;
	assign cst_8_in1_valid = source_4_out1_valid;
	assign source_4_out1_ready = cst_8_in1_ready;

	assign source_5_clk = clk;
	assign source_5_rst = rst;
	assign cst_9_in1_data = source_5_out1_data;
	assign cst_9_in1_valid = source_5_out1_valid;
	assign source_5_out1_ready = cst_9_in1_ready;

	assign source_6_clk = clk;
	assign source_6_rst = rst;
	assign cst_10_in1_data = source_6_out1_data;
	assign cst_10_in1_valid = source_6_out1_valid;
	assign source_6_out1_ready = cst_10_in1_ready;

	assign ret_0_clk = clk;
	assign ret_0_rst = rst;
	assign end_0_in4_data = ret_0_out1_data;
	assign end_0_in4_valid = ret_0_out1_valid;
	assign ret_0_out1_ready = end_0_in4_ready;

	assign end_0_clk = clk;
	assign end_0_rst = rst;
	assign end_out = end_0_out1_data;
	assign end_0_out1_ready = end_ready;
	assign end_valid = end_0_out1_valid;

	assign phiC_12_clk = clk;
	assign phiC_12_rst = rst;
	assign ret_0_in1_data = phiC_12_out1_data;
	assign ret_0_in1_valid = phiC_12_out1_valid;
	assign phiC_12_out1_ready = ret_0_in1_ready;

	assign phi_1_clk = clk;
	assign phi_1_rst = rst;
	assign branch_2_in1_data = phi_1_out1_data;
	assign branch_2_in1_valid = phi_1_out1_valid;
	assign phi_1_out1_ready = branch_2_in1_ready;

	assign brCst_block2_clk = clk;
	assign brCst_block2_rst = rst;
	assign fork_10_in1_data = brCst_block2_out1_data;
	assign fork_10_in1_valid = brCst_block2_out1_valid;
	assign brCst_block2_out1_ready = fork_10_in1_ready;

	assign cst_1_clk = clk;
	assign cst_1_rst = rst;
	assign branch_1_in1_data = cst_1_out1_data;
	assign branch_1_in1_valid = cst_1_out1_valid;
	assign cst_1_out1_ready = branch_1_in1_ready;

	assign branch_1_clk = clk;
	assign branch_1_rst = rst;
	assign phi_3_in2_data = branch_1_out1_data;
	assign phi_3_in2_valid = branch_1_out1_valid;
	assign branch_1_out1_ready = phi_3_in2_ready;
	assign sink_1_in1_data = branch_1_out2_data;
	assign sink_1_in1_valid = branch_1_out2_valid;
	assign branch_1_out2_ready = sink_1_in1_ready;

	assign branch_2_clk = clk;
	assign branch_2_rst = rst;
	assign phi_n1_in1_data = branch_2_out1_data;
	assign phi_n1_in1_valid = branch_2_out1_valid;
	assign branch_2_out1_ready = phi_n1_in1_ready;
	assign sink_2_in1_data = branch_2_out2_data;
	assign sink_2_in1_valid = branch_2_out2_valid;
	assign branch_2_out2_ready = sink_2_in1_ready;

	assign fork_10_clk = clk;
	assign fork_10_rst = rst;
	assign branch_2_in2_data = fork_10_out1_data;
	assign branch_2_in2_valid = fork_10_out1_valid;
	assign fork_10_out1_ready = branch_2_in2_ready;
	assign branch_1_in2_data = fork_10_out2_data;
	assign branch_1_in2_valid = fork_10_out2_valid;
	assign fork_10_out2_ready = branch_1_in2_ready;
	assign branchC_15_in2_data = fork_10_out3_data;
	assign branchC_15_in2_valid = fork_10_out3_valid;
	assign fork_10_out3_ready = branchC_15_in2_ready;

	assign phiC_7_clk = clk;
	assign phiC_7_rst = rst;
	assign forkC_18_in1_data = phiC_7_out1_data;
	assign forkC_18_in1_valid = phiC_7_out1_valid;
	assign phiC_7_out1_ready = forkC_18_in1_ready;
	assign phi_1_in1_data = phiC_7_out2_data;
	assign phi_1_in1_valid = phiC_7_out2_valid;
	assign phiC_7_out2_ready = phi_1_in1_ready;

	assign forkC_18_clk = clk;
	assign forkC_18_rst = rst;
	assign cst_1_in1_data = forkC_18_out1_data;
	assign cst_1_in1_valid = forkC_18_out1_valid;
	assign forkC_18_out1_ready = cst_1_in1_ready;
	assign branchC_15_in1_data = forkC_18_out2_data;
	assign branchC_15_in1_valid = forkC_18_out2_valid;
	assign forkC_18_out2_ready = branchC_15_in1_ready;
	assign brCst_block2_in1_data = forkC_18_out3_data;
	assign brCst_block2_in1_valid = forkC_18_out3_valid;
	assign forkC_18_out3_ready = brCst_block2_in1_ready;

	assign branchC_15_clk = clk;
	assign branchC_15_rst = rst;
	assign phiC_8_in1_data = branchC_15_out1_data;
	assign phiC_8_in1_valid = branchC_15_out1_valid;
	assign branchC_15_out1_ready = phiC_8_in1_ready;
	assign sink_11_in1_data = branchC_15_out2_data;
	assign sink_11_in1_valid = branchC_15_out2_valid;
	assign branchC_15_out2_ready = sink_11_in1_ready;

	assign MC_in_a_clk = clk;
	assign MC_in_a_rst = rst;
	assign in_a_ce0 = in_a_we0;
	assign MC_in_a_in2_valid = 0;
	assign MC_in_a_in2_data = 0;
	assign load_11_in1_data = MC_in_a_out1_data;
	assign load_11_in1_valid = MC_in_a_out1_valid;
	assign MC_in_a_out1_ready = load_11_in1_ready;
	assign end_0_in1_data = MC_in_a_out2_data;
	assign end_0_in1_valid = MC_in_a_out2_valid;
	assign MC_in_a_out2_ready = end_0_in1_ready;

	assign MC_in_b_clk = clk;
	assign MC_in_b_rst = rst;
	assign in_b_ce0 = in_b_we0;
	assign MC_in_b_in2_valid = 0;
	assign MC_in_b_in2_data = 0;
	assign load_16_in1_data = MC_in_b_out1_data;
	assign load_16_in1_valid = MC_in_b_out1_valid;
	assign MC_in_b_out1_ready = load_16_in1_ready;
	assign end_0_in2_data = MC_in_b_out2_data;
	assign end_0_in2_valid = MC_in_b_out2_valid;
	assign MC_in_b_out2_ready = end_0_in2_ready;

	assign MC_out_c_clk = clk;
	assign MC_out_c_rst = rst;
	assign out_c_ce0 = out_c_we0;
	assign end_0_in3_data = MC_out_c_out1_data;
	assign end_0_in3_valid = MC_out_c_out1_valid;
	assign MC_out_c_out1_ready = end_0_in3_ready;

	assign sink_0_clk = clk;
	assign sink_0_rst = rst;

	assign sink_1_clk = clk;
	assign sink_1_rst = rst;

	assign sink_2_clk = clk;
	assign sink_2_rst = rst;

	assign sink_3_clk = clk;
	assign sink_3_rst = rst;

	assign sink_4_clk = clk;
	assign sink_4_rst = rst;

	assign sink_5_clk = clk;
	assign sink_5_rst = rst;

	assign sink_6_clk = clk;
	assign sink_6_rst = rst;

	assign sink_7_clk = clk;
	assign sink_7_rst = rst;

	assign sink_8_clk = clk;
	assign sink_8_rst = rst;

	assign sink_9_clk = clk;
	assign sink_9_rst = rst;

	assign sink_10_clk = clk;
	assign sink_10_rst = rst;

	assign sink_11_clk = clk;
	assign sink_11_rst = rst;

	assign sink_12_clk = clk;
	assign sink_12_rst = rst;

	assign Buffer_100_clk = clk;
	assign Buffer_100_rst = rst;
	assign phi_5_in3_data = Buffer_100_out1_data;
	assign phi_5_in3_valid = Buffer_100_out1_valid;
	assign Buffer_100_out1_ready = phi_5_in3_ready;

	assign Buffer_101_clk = clk;
	assign Buffer_101_rst = rst;
	assign phi_6_in3_data = Buffer_101_out1_data;
	assign phi_6_in3_valid = Buffer_101_out1_valid;
	assign Buffer_101_out1_ready = phi_6_in3_ready;

	assign Buffer_102_clk = clk;
	assign Buffer_102_rst = rst;
	assign phi_n5_in2_data = Buffer_102_out1_data;
	assign phi_n5_in2_valid = Buffer_102_out1_valid;
	assign Buffer_102_out1_ready = phi_n5_in2_ready;

	assign Buffer_103_clk = clk;
	assign Buffer_103_rst = rst;
	assign phi_n6_in2_data = Buffer_103_out1_data;
	assign phi_n6_in2_valid = Buffer_103_out1_valid;
	assign Buffer_103_out1_ready = phi_n6_in2_ready;

	assign Buffer_104_clk = clk;
	assign Buffer_104_rst = rst;
	assign phiC_9_in2_data = Buffer_104_out1_data;
	assign phiC_9_in2_valid = Buffer_104_out1_valid;
	assign Buffer_104_out1_ready = phiC_9_in2_ready;

	assign Buffer_105_clk = clk;
	assign Buffer_105_rst = rst;
	assign phi_3_in3_data = Buffer_105_out1_data;
	assign phi_3_in3_valid = Buffer_105_out1_valid;
	assign Buffer_105_out1_ready = phi_3_in3_ready;

	assign Buffer_106_clk = clk;
	assign Buffer_106_rst = rst;
	assign phi_n1_in2_data = Buffer_106_out1_data;
	assign phi_n1_in2_valid = Buffer_106_out1_valid;
	assign Buffer_106_out1_ready = phi_n1_in2_ready;

	assign Buffer_107_clk = clk;
	assign Buffer_107_rst = rst;
	assign phiC_8_in2_data = Buffer_107_out1_data;
	assign phiC_8_in2_valid = Buffer_107_out1_valid;
	assign Buffer_107_out1_ready = phiC_8_in2_ready;

	assign Buffer_108_clk = clk;
	assign Buffer_108_rst = rst;
	assign phi_1_in3_data = Buffer_108_out1_data;
	assign phi_1_in3_valid = Buffer_108_out1_valid;
	assign Buffer_108_out1_ready = phi_1_in3_ready;

	assign Buffer_109_clk = clk;
	assign Buffer_109_rst = rst;
	assign phiC_7_in2_data = Buffer_109_out1_data;
	assign phiC_7_in2_valid = Buffer_109_out1_valid;
	assign Buffer_109_out1_ready = phiC_7_in2_ready;

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block1
		(.clk(brCst_block1_clk), .rst(brCst_block1_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block1_in1_valid}), .ready_in_bus({brCst_block1_in1_ready}), 
		.data_out_bus({brCst_block1_out1_data}), .valid_out_bus({brCst_block1_out1_valid}), .ready_out_bus({brCst_block1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_0
		(.clk(cst_0_clk), .rst(cst_0_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_0_in1_valid}), .ready_in_bus({cst_0_in1_ready}), 
		.data_out_bus({cst_0_out1_data}), .valid_out_bus({cst_0_out1_valid}), .ready_out_bus({cst_0_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_0
		(.clk(branch_0_clk), .rst(branch_0_rst),
		.data_in_bus({{branch_0_in2_data}, branch_0_in1_data}), .valid_in_bus({branch_0_in2_valid, branch_0_in1_valid}), .ready_in_bus({branch_0_in2_ready, branch_0_in1_ready}), 
		.data_out_bus({branch_0_out2_data, branch_0_out1_data}), .valid_out_bus({branch_0_out2_valid, branch_0_out1_valid}), .ready_out_bus({branch_0_out2_ready, branch_0_out1_ready}));

	start_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) start_node_start_0
		(.clk(start_0_clk), .rst(start_0_rst),
		.data_in_bus({start_0_in1_data}), .valid_in_bus({start_0_in1_valid}), .ready_in_bus({start_0_in1_ready}), 
		.data_out_bus({start_0_out1_data}), .valid_out_bus({start_0_out1_valid}), .ready_out_bus({start_0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_16
		(.clk(forkC_16_clk), .rst(forkC_16_rst),
		.data_in_bus({forkC_16_in1_data}), .valid_in_bus({forkC_16_in1_valid}), .ready_in_bus({forkC_16_in1_ready}), 
		.data_out_bus({forkC_16_out3_data, forkC_16_out2_data, forkC_16_out1_data}), .valid_out_bus({forkC_16_out3_valid, forkC_16_out2_valid, forkC_16_out1_valid}), .ready_out_bus({forkC_16_out3_ready, forkC_16_out2_ready, forkC_16_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_14
		(.clk(branchC_14_clk), .rst(branchC_14_rst),
		.data_in_bus({{branchC_14_in2_data}, branchC_14_in1_data}), .valid_in_bus({branchC_14_in2_valid, branchC_14_in1_valid}), .ready_in_bus({branchC_14_in2_ready, branchC_14_in1_ready}), 
		.data_out_bus({branchC_14_out2_data, branchC_14_out1_data}), .valid_out_bus({branchC_14_out2_valid, branchC_14_out1_valid}), .ready_out_bus({branchC_14_out2_ready, branchC_14_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_17
		(.clk(fork_17_clk), .rst(fork_17_rst),
		.data_in_bus({fork_17_in1_data}), .valid_in_bus({fork_17_in1_valid}), .ready_in_bus({fork_17_in1_ready}), 
		.data_out_bus({fork_17_out2_data, fork_17_out1_data}), .valid_out_bus({fork_17_out2_valid, fork_17_out1_valid}), .ready_out_bus({fork_17_out2_ready, fork_17_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_3
		(.clk(phi_3_clk), .rst(phi_3_rst),
		.data_in_bus({{5'b0, phi_3_in1_data}, phi_3_in3_data, phi_3_in2_data}), .valid_in_bus({phi_3_in1_valid, phi_3_in3_valid, phi_3_in2_valid}), .ready_in_bus({phi_3_in1_ready, phi_3_in3_ready, phi_3_in2_ready}), 
		.data_out_bus({phi_3_out1_data}), .valid_out_bus({phi_3_out1_valid}), .ready_out_bus({phi_3_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block3
		(.clk(brCst_block3_clk), .rst(brCst_block3_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block3_in1_valid}), .ready_in_bus({brCst_block3_in1_ready}), 
		.data_out_bus({brCst_block3_out1_data}), .valid_out_bus({brCst_block3_out1_valid}), .ready_out_bus({brCst_block3_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_2
		(.clk(cst_2_clk), .rst(cst_2_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_2_in1_valid}), .ready_in_bus({cst_2_in1_ready}), 
		.data_out_bus({cst_2_out1_data}), .valid_out_bus({cst_2_out1_valid}), .ready_out_bus({cst_2_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_3
		(.clk(cst_3_clk), .rst(cst_3_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_3_in1_valid}), .ready_in_bus({cst_3_in1_ready}), 
		.data_out_bus({cst_3_out1_data}), .valid_out_bus({cst_3_out1_valid}), .ready_out_bus({cst_3_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n1
		(.clk(phi_n1_clk), .rst(phi_n1_rst),
		.data_in_bus({phi_n1_in2_data, phi_n1_in1_data}), .valid_in_bus({phi_n1_in2_valid, phi_n1_in1_valid}), .ready_in_bus({phi_n1_in2_ready, phi_n1_in1_ready}), 
		.data_out_bus({phi_n1_out1_data}), .valid_out_bus({phi_n1_out1_valid}), .ready_out_bus({phi_n1_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_3
		(.clk(branch_3_clk), .rst(branch_3_rst),
		.data_in_bus({{branch_3_in2_data}, branch_3_in1_data}), .valid_in_bus({branch_3_in2_valid, branch_3_in1_valid}), .ready_in_bus({branch_3_in2_ready, branch_3_in1_ready}), 
		.data_out_bus({branch_3_out2_data, branch_3_out1_data}), .valid_out_bus({branch_3_out2_valid, branch_3_out1_valid}), .ready_out_bus({branch_3_out2_ready, branch_3_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_4
		(.clk(branch_4_clk), .rst(branch_4_rst),
		.data_in_bus({{branch_4_in2_data}, branch_4_in1_data}), .valid_in_bus({branch_4_in2_valid, branch_4_in1_valid}), .ready_in_bus({branch_4_in2_ready, branch_4_in1_ready}), 
		.data_out_bus({branch_4_out2_data, branch_4_out1_data}), .valid_out_bus({branch_4_out2_valid, branch_4_out1_valid}), .ready_out_bus({branch_4_out2_ready, branch_4_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_5
		(.clk(branch_5_clk), .rst(branch_5_rst),
		.data_in_bus({{5'b0, branch_5_in2_data}, branch_5_in1_data}), .valid_in_bus({branch_5_in2_valid, branch_5_in1_valid}), .ready_in_bus({branch_5_in2_ready, branch_5_in1_ready}), 
		.data_out_bus({branch_5_out2_data, branch_5_out1_data}), .valid_out_bus({branch_5_out2_valid, branch_5_out1_valid}), .ready_out_bus({branch_5_out2_ready, branch_5_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_6
		(.clk(branch_6_clk), .rst(branch_6_rst),
		.data_in_bus({{5'b0, branch_6_in2_data}, branch_6_in1_data}), .valid_in_bus({branch_6_in2_valid, branch_6_in1_valid}), .ready_in_bus({branch_6_in2_ready, branch_6_in1_ready}), 
		.data_out_bus({branch_6_out2_data, branch_6_out1_data}), .valid_out_bus({branch_6_out2_valid, branch_6_out1_valid}), .ready_out_bus({branch_6_out2_ready, branch_6_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_11
		(.clk(fork_11_clk), .rst(fork_11_rst),
		.data_in_bus({fork_11_in1_data}), .valid_in_bus({fork_11_in1_valid}), .ready_in_bus({fork_11_in1_ready}), 
		.data_out_bus({fork_11_out5_data, fork_11_out4_data, fork_11_out3_data, fork_11_out2_data, fork_11_out1_data}), .valid_out_bus({fork_11_out5_valid, fork_11_out4_valid, fork_11_out3_valid, fork_11_out2_valid, fork_11_out1_valid}), .ready_out_bus({fork_11_out5_ready, fork_11_out4_ready, fork_11_out3_ready, fork_11_out2_ready, fork_11_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_8
		(.clk(phiC_8_clk), .rst(phiC_8_rst),
		.data_in_bus({phiC_8_in2_data, phiC_8_in1_data}), .valid_in_bus({phiC_8_in2_valid, phiC_8_in1_valid}), .ready_in_bus({phiC_8_in2_ready, phiC_8_in1_ready}), 
		.data_out_bus({phiC_8_out2_data, phiC_8_out1_data}), .valid_out_bus({phiC_8_out2_valid, phiC_8_out1_valid}), .ready_out_bus({phiC_8_out2_ready, phiC_8_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_19
		(.clk(forkC_19_clk), .rst(forkC_19_rst),
		.data_in_bus({forkC_19_in1_data}), .valid_in_bus({forkC_19_in1_valid}), .ready_in_bus({forkC_19_in1_ready}), 
		.data_out_bus({forkC_19_out4_data, forkC_19_out3_data, forkC_19_out2_data, forkC_19_out1_data}), .valid_out_bus({forkC_19_out4_valid, forkC_19_out3_valid, forkC_19_out2_valid, forkC_19_out1_valid}), .ready_out_bus({forkC_19_out4_ready, forkC_19_out3_ready, forkC_19_out2_ready, forkC_19_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_16
		(.clk(branchC_16_clk), .rst(branchC_16_rst),
		.data_in_bus({{branchC_16_in2_data}, branchC_16_in1_data}), .valid_in_bus({branchC_16_in2_valid, branchC_16_in1_valid}), .ready_in_bus({branchC_16_in2_ready, branchC_16_in1_ready}), 
		.data_out_bus({branchC_16_out2_data, branchC_16_out1_data}), .valid_out_bus({branchC_16_out2_valid, branchC_16_out1_valid}), .ready_out_bus({branchC_16_out2_ready, branchC_16_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_11
		(.clk(cst_11_clk), .rst(cst_11_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_11_in1_valid}), .ready_in_bus({cst_11_in1_ready}), 
		.data_out_bus({cst_11_out1_data}), .valid_out_bus({cst_11_out1_valid}), .ready_out_bus({cst_11_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_29
		(.clk(add_29_clk), .rst(add_29_rst),
		.data_in_bus({add_29_in2_data, add_29_in1_data}), .valid_in_bus({add_29_in2_valid, add_29_in1_valid}), .ready_in_bus({add_29_in2_ready, add_29_in1_ready}), 
		.data_out_bus({add_29_out1_data}), .valid_out_bus({add_29_out1_valid}), .ready_out_bus({add_29_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_12
		(.clk(cst_12_clk), .rst(cst_12_rst),
		.data_in_bus({6'd32}), .valid_in_bus({cst_12_in1_valid}), .ready_in_bus({cst_12_in1_ready}), 
		.data_out_bus({cst_12_out1_data}), .valid_out_bus({cst_12_out1_valid}), .ready_out_bus({cst_12_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_30
		(.clk(icmp_30_clk), .rst(icmp_30_rst),
		.data_in_bus({icmp_30_in2_data, icmp_30_in1_data}), .valid_in_bus({icmp_30_in2_valid, icmp_30_in1_valid}), .ready_in_bus({icmp_30_in2_ready, icmp_30_in1_ready}), 
		.data_out_bus({icmp_30_out1_data}), .valid_out_bus({icmp_30_out1_valid}), .ready_out_bus({icmp_30_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n0
		(.clk(phi_n0_clk), .rst(phi_n0_rst),
		.data_in_bus({phi_n0_in1_data}), .valid_in_bus({phi_n0_in1_valid}), .ready_in_bus({phi_n0_in1_ready}), 
		.data_out_bus({phi_n0_out1_data}), .valid_out_bus({phi_n0_out1_valid}), .ready_out_bus({phi_n0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_4
		(.clk(fork_4_clk), .rst(fork_4_rst),
		.data_in_bus({fork_4_in1_data}), .valid_in_bus({fork_4_in1_valid}), .ready_in_bus({fork_4_in1_ready}), 
		.data_out_bus({fork_4_out2_data, fork_4_out1_data}), .valid_out_bus({fork_4_out2_valid, fork_4_out1_valid}), .ready_out_bus({fork_4_out2_ready, fork_4_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_13
		(.clk(branch_13_clk), .rst(branch_13_rst),
		.data_in_bus({{5'b0, branch_13_in2_data}, branch_13_in1_data}), .valid_in_bus({branch_13_in2_valid, branch_13_in1_valid}), .ready_in_bus({branch_13_in2_ready, branch_13_in1_ready}), 
		.data_out_bus({branch_13_out2_data, branch_13_out1_data}), .valid_out_bus({branch_13_out2_valid, branch_13_out1_valid}), .ready_out_bus({branch_13_out2_ready, branch_13_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_11
		(.clk(phiC_11_clk), .rst(phiC_11_rst),
		.data_in_bus({phiC_11_in1_data}), .valid_in_bus({phiC_11_in1_valid}), .ready_in_bus({phiC_11_in1_ready}), 
		.data_out_bus({phiC_11_out1_data}), .valid_out_bus({phiC_11_out1_valid}), .ready_out_bus({phiC_11_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_19
		(.clk(branchC_19_clk), .rst(branchC_19_rst),
		.data_in_bus({{branchC_19_in2_data}, branchC_19_in1_data}), .valid_in_bus({branchC_19_in2_valid, branchC_19_in1_valid}), .ready_in_bus({branchC_19_in2_ready, branchC_19_in1_ready}), 
		.data_out_bus({branchC_19_out2_data, branchC_19_out1_data}), .valid_out_bus({branchC_19_out2_valid, branchC_19_out1_valid}), .ready_out_bus({branchC_19_out2_ready, branchC_19_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_23
		(.clk(fork_23_clk), .rst(fork_23_rst),
		.data_in_bus({fork_23_in1_data}), .valid_in_bus({fork_23_in1_valid}), .ready_in_bus({fork_23_in1_ready}), 
		.data_out_bus({fork_23_out2_data, fork_23_out1_data}), .valid_out_bus({fork_23_out2_valid, fork_23_out1_valid}), .ready_out_bus({fork_23_out2_ready, fork_23_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_7
		(.clk(source_7_clk), .rst(source_7_rst),
		.data_out_bus({source_7_out1_data}), .valid_out_bus({source_7_out1_valid}), .ready_out_bus({source_7_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_8
		(.clk(source_8_clk), .rst(source_8_rst),
		.data_out_bus({source_8_out1_data}), .valid_out_bus({source_8_out1_valid}), .ready_out_bus({source_8_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_5
		(.clk(phi_5_clk), .rst(phi_5_rst),
		.data_in_bus({{31'b0, phi_5_in1_data}, phi_5_in3_data, phi_5_in2_data}), .valid_in_bus({phi_5_in1_valid, phi_5_in3_valid, phi_5_in2_valid}), .ready_in_bus({phi_5_in1_ready, phi_5_in3_ready, phi_5_in2_ready}), 
		.data_out_bus({phi_5_out1_data}), .valid_out_bus({phi_5_out1_valid}), .ready_out_bus({phi_5_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_6
		(.clk(phi_6_clk), .rst(phi_6_rst),
		.data_in_bus({{5'b0, phi_6_in1_data}, phi_6_in3_data, phi_6_in2_data}), .valid_in_bus({phi_6_in1_valid, phi_6_in3_valid, phi_6_in2_valid}), .ready_in_bus({phi_6_in1_ready, phi_6_in3_ready, phi_6_in2_ready}), 
		.data_out_bus({phi_6_out1_data}), .valid_out_bus({phi_6_out1_valid}), .ready_out_bus({phi_6_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_4
		(.clk(cst_4_clk), .rst(cst_4_rst),
		.data_in_bus({3'd5}), .valid_in_bus({cst_4_in1_valid}), .ready_in_bus({cst_4_in1_ready}), 
		.data_out_bus({cst_4_out1_data}), .valid_out_bus({cst_4_out1_valid}), .ready_out_bus({cst_4_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(11), .DATA_OUT_SIZE(11)) shl_op_shl_7
		(.clk(shl_7_clk), .rst(shl_7_rst),
		.data_in_bus({shl_7_in2_data, shl_7_in1_data}), .valid_in_bus({shl_7_in2_valid, shl_7_in1_valid}), .ready_in_bus({shl_7_in2_ready, shl_7_in1_ready}), 
		.data_out_bus({shl_7_out1_data}), .valid_out_bus({shl_7_out1_valid}), .ready_out_bus({shl_7_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(12), .DATA_OUT_SIZE(12)) add_op_add_8
		(.clk(add_8_clk), .rst(add_8_rst),
		.data_in_bus({add_8_in2_data, add_8_in1_data}), .valid_in_bus({add_8_in2_valid, add_8_in1_valid}), .ready_in_bus({add_8_in2_ready, add_8_in1_ready}), 
		.data_out_bus({add_8_out1_data}), .valid_out_bus({add_8_out1_valid}), .ready_out_bus({add_8_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(12), .DATA_SIZE(32)) mc_load_op_load_11
		(.clk(load_11_clk), .rst(load_11_rst),
		.data_in_bus({load_11_in1_data}), .address_in_bus({load_11_in2_data}), .valid_in_bus({load_11_in2_valid, load_11_in1_valid}), .ready_in_bus({load_11_in2_ready, load_11_in1_ready}), 
		.data_out_bus({load_11_out1_data}), .address_out_bus({load_11_out2_data}), .valid_out_bus({load_11_out2_valid, load_11_out1_valid}), .ready_out_bus({load_11_out2_ready, load_11_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_5
		(.clk(cst_5_clk), .rst(cst_5_rst),
		.data_in_bus({3'd5}), .valid_in_bus({cst_5_in1_valid}), .ready_in_bus({cst_5_in1_ready}), 
		.data_out_bus({cst_5_out1_data}), .valid_out_bus({cst_5_out1_valid}), .ready_out_bus({cst_5_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(11), .DATA_OUT_SIZE(11)) shl_op_shl_12
		(.clk(shl_12_clk), .rst(shl_12_rst),
		.data_in_bus({shl_12_in2_data, shl_12_in1_data}), .valid_in_bus({shl_12_in2_valid, shl_12_in1_valid}), .ready_in_bus({shl_12_in2_ready, shl_12_in1_ready}), 
		.data_out_bus({shl_12_out1_data}), .valid_out_bus({shl_12_out1_valid}), .ready_out_bus({shl_12_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(12), .DATA_OUT_SIZE(12)) add_op_add_13
		(.clk(add_13_clk), .rst(add_13_rst),
		.data_in_bus({add_13_in2_data, add_13_in1_data}), .valid_in_bus({add_13_in2_valid, add_13_in1_valid}), .ready_in_bus({add_13_in2_ready, add_13_in1_ready}), 
		.data_out_bus({add_13_out1_data}), .valid_out_bus({add_13_out1_valid}), .ready_out_bus({add_13_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(12), .DATA_SIZE(32)) mc_load_op_load_16
		(.clk(load_16_clk), .rst(load_16_rst),
		.data_in_bus({load_16_in1_data}), .address_in_bus({load_16_in2_data}), .valid_in_bus({load_16_in2_valid, load_16_in1_valid}), .ready_in_bus({load_16_in2_ready, load_16_in1_ready}), 
		.data_out_bus({load_16_out1_data}), .address_out_bus({load_16_out2_data}), .valid_out_bus({load_16_out2_valid, load_16_out1_valid}), .ready_out_bus({load_16_out2_ready, load_16_out1_ready}));

	mul_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(16), .DATA_OUT_SIZE(32)) mul_op_mul_17
		(.clk(mul_17_clk), .rst(mul_17_rst),
		.data_in_bus({mul_17_in2_data, mul_17_in1_data}), .valid_in_bus({mul_17_in2_valid, mul_17_in1_valid}), .ready_in_bus({mul_17_in2_ready, mul_17_in1_ready}), 
		.data_out_bus({mul_17_out1_data}), .valid_out_bus({mul_17_out1_valid}), .ready_out_bus({mul_17_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_18
		(.clk(add_18_clk), .rst(add_18_rst),
		.data_in_bus({add_18_in2_data, add_18_in1_data}), .valid_in_bus({add_18_in2_valid, add_18_in1_valid}), .ready_in_bus({add_18_in2_ready, add_18_in1_ready}), 
		.data_out_bus({add_18_out1_data}), .valid_out_bus({add_18_out1_valid}), .ready_out_bus({add_18_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_6
		(.clk(cst_6_clk), .rst(cst_6_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_6_in1_valid}), .ready_in_bus({cst_6_in1_ready}), 
		.data_out_bus({cst_6_out1_data}), .valid_out_bus({cst_6_out1_valid}), .ready_out_bus({cst_6_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_19
		(.clk(add_19_clk), .rst(add_19_rst),
		.data_in_bus({add_19_in2_data, add_19_in1_data}), .valid_in_bus({add_19_in2_valid, add_19_in1_valid}), .ready_in_bus({add_19_in2_ready, add_19_in1_ready}), 
		.data_out_bus({add_19_out1_data}), .valid_out_bus({add_19_out1_valid}), .ready_out_bus({add_19_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_7
		(.clk(cst_7_clk), .rst(cst_7_rst),
		.data_in_bus({6'd32}), .valid_in_bus({cst_7_in1_valid}), .ready_in_bus({cst_7_in1_ready}), 
		.data_out_bus({cst_7_out1_data}), .valid_out_bus({cst_7_out1_valid}), .ready_out_bus({cst_7_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_20
		(.clk(icmp_20_clk), .rst(icmp_20_rst),
		.data_in_bus({icmp_20_in2_data, icmp_20_in1_data}), .valid_in_bus({icmp_20_in2_valid, icmp_20_in1_valid}), .ready_in_bus({icmp_20_in2_ready, icmp_20_in1_ready}), 
		.data_out_bus({icmp_20_out1_data}), .valid_out_bus({icmp_20_out1_valid}), .ready_out_bus({icmp_20_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n5
		(.clk(phi_n5_clk), .rst(phi_n5_rst),
		.data_in_bus({phi_n5_in2_data, phi_n5_in1_data}), .valid_in_bus({phi_n5_in2_valid, phi_n5_in1_valid}), .ready_in_bus({phi_n5_in2_ready, phi_n5_in1_ready}), 
		.data_out_bus({phi_n5_out1_data}), .valid_out_bus({phi_n5_out1_valid}), .ready_out_bus({phi_n5_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n6
		(.clk(phi_n6_clk), .rst(phi_n6_rst),
		.data_in_bus({phi_n6_in2_data, phi_n6_in1_data}), .valid_in_bus({phi_n6_in2_valid, phi_n6_in1_valid}), .ready_in_bus({phi_n6_in2_ready, phi_n6_in1_ready}), 
		.data_out_bus({phi_n6_out1_data}), .valid_out_bus({phi_n6_out1_valid}), .ready_out_bus({phi_n6_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_0
		(.clk(fork_0_clk), .rst(fork_0_rst),
		.data_in_bus({fork_0_in1_data}), .valid_in_bus({fork_0_in1_valid}), .ready_in_bus({fork_0_in1_ready}), 
		.data_out_bus({fork_0_out3_data, fork_0_out2_data, fork_0_out1_data}), .valid_out_bus({fork_0_out3_valid, fork_0_out2_valid, fork_0_out1_valid}), .ready_out_bus({fork_0_out3_ready, fork_0_out2_ready, fork_0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_2
		(.clk(fork_2_clk), .rst(fork_2_rst),
		.data_in_bus({fork_2_in1_data}), .valid_in_bus({fork_2_in1_valid}), .ready_in_bus({fork_2_in1_ready}), 
		.data_out_bus({fork_2_out2_data, fork_2_out1_data}), .valid_out_bus({fork_2_out2_valid, fork_2_out1_valid}), .ready_out_bus({fork_2_out2_ready, fork_2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_7
		(.clk(fork_7_clk), .rst(fork_7_rst),
		.data_in_bus({fork_7_in1_data}), .valid_in_bus({fork_7_in1_valid}), .ready_in_bus({fork_7_in1_ready}), 
		.data_out_bus({fork_7_out2_data, fork_7_out1_data}), .valid_out_bus({fork_7_out2_valid, fork_7_out1_valid}), .ready_out_bus({fork_7_out2_ready, fork_7_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_8
		(.clk(fork_8_clk), .rst(fork_8_rst),
		.data_in_bus({fork_8_in1_data}), .valid_in_bus({fork_8_in1_valid}), .ready_in_bus({fork_8_in1_ready}), 
		.data_out_bus({fork_8_out2_data, fork_8_out1_data}), .valid_out_bus({fork_8_out2_valid, fork_8_out1_valid}), .ready_out_bus({fork_8_out2_ready, fork_8_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_7
		(.clk(branch_7_clk), .rst(branch_7_rst),
		.data_in_bus({{31'b0, branch_7_in2_data}, branch_7_in1_data}), .valid_in_bus({branch_7_in2_valid, branch_7_in1_valid}), .ready_in_bus({branch_7_in2_ready, branch_7_in1_ready}), 
		.data_out_bus({branch_7_out2_data, branch_7_out1_data}), .valid_out_bus({branch_7_out2_valid, branch_7_out1_valid}), .ready_out_bus({branch_7_out2_ready, branch_7_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_8
		(.clk(branch_8_clk), .rst(branch_8_rst),
		.data_in_bus({{5'b0, branch_8_in2_data}, branch_8_in1_data}), .valid_in_bus({branch_8_in2_valid, branch_8_in1_valid}), .ready_in_bus({branch_8_in2_ready, branch_8_in1_ready}), 
		.data_out_bus({branch_8_out2_data, branch_8_out1_data}), .valid_out_bus({branch_8_out2_valid, branch_8_out1_valid}), .ready_out_bus({branch_8_out2_ready, branch_8_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_9
		(.clk(branch_9_clk), .rst(branch_9_rst),
		.data_in_bus({{5'b0, branch_9_in2_data}, branch_9_in1_data}), .valid_in_bus({branch_9_in2_valid, branch_9_in1_valid}), .ready_in_bus({branch_9_in2_ready, branch_9_in1_ready}), 
		.data_out_bus({branch_9_out2_data, branch_9_out1_data}), .valid_out_bus({branch_9_out2_valid, branch_9_out1_valid}), .ready_out_bus({branch_9_out2_ready, branch_9_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_10
		(.clk(branch_10_clk), .rst(branch_10_rst),
		.data_in_bus({{5'b0, branch_10_in2_data}, branch_10_in1_data}), .valid_in_bus({branch_10_in2_valid, branch_10_in1_valid}), .ready_in_bus({branch_10_in2_ready, branch_10_in1_ready}), 
		.data_out_bus({branch_10_out2_data, branch_10_out1_data}), .valid_out_bus({branch_10_out2_valid, branch_10_out1_valid}), .ready_out_bus({branch_10_out2_ready, branch_10_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_12
		(.clk(fork_12_clk), .rst(fork_12_rst),
		.data_in_bus({fork_12_in1_data}), .valid_in_bus({fork_12_in1_valid}), .ready_in_bus({fork_12_in1_ready}), 
		.data_out_bus({fork_12_out5_data, fork_12_out4_data, fork_12_out3_data, fork_12_out2_data, fork_12_out1_data}), .valid_out_bus({fork_12_out5_valid, fork_12_out4_valid, fork_12_out3_valid, fork_12_out2_valid, fork_12_out1_valid}), .ready_out_bus({fork_12_out5_ready, fork_12_out4_ready, fork_12_out3_ready, fork_12_out2_ready, fork_12_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_9
		(.clk(phiC_9_clk), .rst(phiC_9_rst),
		.data_in_bus({phiC_9_in2_data, phiC_9_in1_data}), .valid_in_bus({phiC_9_in2_valid, phiC_9_in1_valid}), .ready_in_bus({phiC_9_in2_ready, phiC_9_in1_ready}), 
		.data_out_bus({phiC_9_out2_data, phiC_9_out1_data}), .valid_out_bus({phiC_9_out2_valid, phiC_9_out1_valid}), .ready_out_bus({phiC_9_out2_ready, phiC_9_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_17
		(.clk(branchC_17_clk), .rst(branchC_17_rst),
		.data_in_bus({{branchC_17_in2_data}, branchC_17_in1_data}), .valid_in_bus({branchC_17_in2_valid, branchC_17_in1_valid}), .ready_in_bus({branchC_17_in2_ready, branchC_17_in1_ready}), 
		.data_out_bus({branchC_17_out2_data, branchC_17_out1_data}), .valid_out_bus({branchC_17_out2_valid, branchC_17_out1_valid}), .ready_out_bus({branchC_17_out2_ready, branchC_17_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_0
		(.clk(source_0_clk), .rst(source_0_rst),
		.data_out_bus({source_0_out1_data}), .valid_out_bus({source_0_out1_valid}), .ready_out_bus({source_0_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_1
		(.clk(source_1_clk), .rst(source_1_rst),
		.data_out_bus({source_1_out1_data}), .valid_out_bus({source_1_out1_valid}), .ready_out_bus({source_1_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_2
		(.clk(source_2_clk), .rst(source_2_rst),
		.data_out_bus({source_2_out1_data}), .valid_out_bus({source_2_out1_valid}), .ready_out_bus({source_2_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_3
		(.clk(source_3_clk), .rst(source_3_rst),
		.data_out_bus({source_3_out1_data}), .valid_out_bus({source_3_out1_valid}), .ready_out_bus({source_3_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_27
		(.clk(fork_27_clk), .rst(fork_27_rst),
		.data_in_bus({fork_27_in1_data}), .valid_in_bus({fork_27_in1_valid}), .ready_in_bus({fork_27_in1_ready}), 
		.data_out_bus({fork_27_out2_data, fork_27_out1_data}), .valid_out_bus({fork_27_out2_valid, fork_27_out1_valid}), .ready_out_bus({fork_27_out2_ready, fork_27_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_8
		(.clk(cst_8_clk), .rst(cst_8_rst),
		.data_in_bus({3'd5}), .valid_in_bus({cst_8_in1_valid}), .ready_in_bus({cst_8_in1_ready}), 
		.data_out_bus({cst_8_out1_data}), .valid_out_bus({cst_8_out1_valid}), .ready_out_bus({cst_8_out1_ready}));

	shl_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(11), .DATA_OUT_SIZE(11)) shl_op_shl_22
		(.clk(shl_22_clk), .rst(shl_22_rst),
		.data_in_bus({shl_22_in2_data, shl_22_in1_data}), .valid_in_bus({shl_22_in2_valid, shl_22_in1_valid}), .ready_in_bus({shl_22_in2_ready, shl_22_in1_ready}), 
		.data_out_bus({shl_22_out1_data}), .valid_out_bus({shl_22_out1_valid}), .ready_out_bus({shl_22_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(12), .DATA_OUT_SIZE(12)) add_op_add_23
		(.clk(add_23_clk), .rst(add_23_rst),
		.data_in_bus({add_23_in2_data, add_23_in1_data}), .valid_in_bus({add_23_in2_valid, add_23_in1_valid}), .ready_in_bus({add_23_in2_ready, add_23_in1_ready}), 
		.data_out_bus({add_23_out1_data}), .valid_out_bus({add_23_out1_valid}), .ready_out_bus({add_23_out1_ready}));

	mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(12), .DATA_SIZE(32)) mc_store_op_store_0
		(.clk(store_0_clk), .rst(store_0_rst),
		.data_in_bus({store_0_in1_data}), .address_in_bus({store_0_in2_data}), .valid_in_bus({store_0_in2_valid, store_0_in1_valid}), .ready_in_bus({store_0_in2_ready, store_0_in1_ready}), 
		.data_out_bus({store_0_out1_data}), .address_out_bus({store_0_out2_data}), .valid_out_bus({store_0_out2_valid, store_0_out1_valid}), .ready_out_bus({store_0_out2_ready, store_0_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_9
		(.clk(cst_9_clk), .rst(cst_9_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_9_in1_valid}), .ready_in_bus({cst_9_in1_ready}), 
		.data_out_bus({cst_9_out1_data}), .valid_out_bus({cst_9_out1_valid}), .ready_out_bus({cst_9_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) add_op_add_26
		(.clk(add_26_clk), .rst(add_26_rst),
		.data_in_bus({add_26_in2_data, add_26_in1_data}), .valid_in_bus({add_26_in2_valid, add_26_in1_valid}), .ready_in_bus({add_26_in2_ready, add_26_in1_ready}), 
		.data_out_bus({add_26_out1_data}), .valid_out_bus({add_26_out1_valid}), .ready_out_bus({add_26_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) const_node_cst_10
		(.clk(cst_10_clk), .rst(cst_10_rst),
		.data_in_bus({6'd32}), .valid_in_bus({cst_10_in1_valid}), .ready_in_bus({cst_10_in1_ready}), 
		.data_out_bus({cst_10_out1_data}), .valid_out_bus({cst_10_out1_valid}), .ready_out_bus({cst_10_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_27
		(.clk(icmp_27_clk), .rst(icmp_27_rst),
		.data_in_bus({icmp_27_in2_data, icmp_27_in1_data}), .valid_in_bus({icmp_27_in2_valid, icmp_27_in1_valid}), .ready_in_bus({icmp_27_in2_ready, icmp_27_in1_ready}), 
		.data_out_bus({icmp_27_out1_data}), .valid_out_bus({icmp_27_out1_valid}), .ready_out_bus({icmp_27_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n2
		(.clk(phi_n2_clk), .rst(phi_n2_rst),
		.data_in_bus({phi_n2_in1_data}), .valid_in_bus({phi_n2_in1_valid}), .ready_in_bus({phi_n2_in1_ready}), 
		.data_out_bus({phi_n2_out1_data}), .valid_out_bus({phi_n2_out1_valid}), .ready_out_bus({phi_n2_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) merge_node_phi_n3
		(.clk(phi_n3_clk), .rst(phi_n3_rst),
		.data_in_bus({phi_n3_in1_data}), .valid_in_bus({phi_n3_in1_valid}), .ready_in_bus({phi_n3_in1_ready}), 
		.data_out_bus({phi_n3_out1_data}), .valid_out_bus({phi_n3_out1_valid}), .ready_out_bus({phi_n3_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n4
		(.clk(phi_n4_clk), .rst(phi_n4_rst),
		.data_in_bus({phi_n4_in1_data}), .valid_in_bus({phi_n4_in1_valid}), .ready_in_bus({phi_n4_in1_ready}), 
		.data_out_bus({phi_n4_out1_data}), .valid_out_bus({phi_n4_out1_valid}), .ready_out_bus({phi_n4_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_3
		(.clk(fork_3_clk), .rst(fork_3_rst),
		.data_in_bus({fork_3_in1_data}), .valid_in_bus({fork_3_in1_valid}), .ready_in_bus({fork_3_in1_ready}), 
		.data_out_bus({fork_3_out2_data, fork_3_out1_data}), .valid_out_bus({fork_3_out2_valid, fork_3_out1_valid}), .ready_out_bus({fork_3_out2_ready, fork_3_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_5
		(.clk(fork_5_clk), .rst(fork_5_rst),
		.data_in_bus({fork_5_in1_data}), .valid_in_bus({fork_5_in1_valid}), .ready_in_bus({fork_5_in1_ready}), 
		.data_out_bus({fork_5_out2_data, fork_5_out1_data}), .valid_out_bus({fork_5_out2_valid, fork_5_out1_valid}), .ready_out_bus({fork_5_out2_ready, fork_5_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) fork_node_fork_6
		(.clk(fork_6_clk), .rst(fork_6_rst),
		.data_in_bus({fork_6_in1_data}), .valid_in_bus({fork_6_in1_valid}), .ready_in_bus({fork_6_in1_ready}), 
		.data_out_bus({fork_6_out2_data, fork_6_out1_data}), .valid_out_bus({fork_6_out2_valid, fork_6_out1_valid}), .ready_out_bus({fork_6_out2_ready, fork_6_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_11
		(.clk(branch_11_clk), .rst(branch_11_rst),
		.data_in_bus({{5'b0, branch_11_in2_data}, branch_11_in1_data}), .valid_in_bus({branch_11_in2_valid, branch_11_in1_valid}), .ready_in_bus({branch_11_in2_ready, branch_11_in1_ready}), 
		.data_out_bus({branch_11_out2_data, branch_11_out1_data}), .valid_out_bus({branch_11_out2_valid, branch_11_out1_valid}), .ready_out_bus({branch_11_out2_ready, branch_11_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_12
		(.clk(branch_12_clk), .rst(branch_12_rst),
		.data_in_bus({{5'b0, branch_12_in2_data}, branch_12_in1_data}), .valid_in_bus({branch_12_in2_valid, branch_12_in1_valid}), .ready_in_bus({branch_12_in2_ready, branch_12_in1_ready}), 
		.data_out_bus({branch_12_out2_data, branch_12_out1_data}), .valid_out_bus({branch_12_out2_valid, branch_12_out1_valid}), .ready_out_bus({branch_12_out2_ready, branch_12_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_13
		(.clk(fork_13_clk), .rst(fork_13_rst),
		.data_in_bus({fork_13_in1_data}), .valid_in_bus({fork_13_in1_valid}), .ready_in_bus({fork_13_in1_ready}), 
		.data_out_bus({fork_13_out3_data, fork_13_out2_data, fork_13_out1_data}), .valid_out_bus({fork_13_out3_valid, fork_13_out2_valid, fork_13_out1_valid}), .ready_out_bus({fork_13_out3_ready, fork_13_out2_ready, fork_13_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_13
		(.clk(cst_13_clk), .rst(cst_13_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_13_in1_valid}), .ready_in_bus({cst_13_in1_ready}), 
		.data_out_bus({cst_13_out1_data}), .valid_out_bus({cst_13_out1_valid}), .ready_out_bus({cst_13_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_10
		(.clk(phiC_10_clk), .rst(phiC_10_rst),
		.data_in_bus({phiC_10_in1_data}), .valid_in_bus({phiC_10_in1_valid}), .ready_in_bus({phiC_10_in1_ready}), 
		.data_out_bus({phiC_10_out1_data}), .valid_out_bus({phiC_10_out1_valid}), .ready_out_bus({phiC_10_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_21
		(.clk(forkC_21_clk), .rst(forkC_21_rst),
		.data_in_bus({forkC_21_in1_data}), .valid_in_bus({forkC_21_in1_valid}), .ready_in_bus({forkC_21_in1_ready}), 
		.data_out_bus({forkC_21_out2_data, forkC_21_out1_data}), .valid_out_bus({forkC_21_out2_valid, forkC_21_out1_valid}), .ready_out_bus({forkC_21_out2_ready, forkC_21_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_18
		(.clk(branchC_18_clk), .rst(branchC_18_rst),
		.data_in_bus({{branchC_18_in2_data}, branchC_18_in1_data}), .valid_in_bus({branchC_18_in2_valid, branchC_18_in1_valid}), .ready_in_bus({branchC_18_in2_ready, branchC_18_in1_ready}), 
		.data_out_bus({branchC_18_out2_data, branchC_18_out1_data}), .valid_out_bus({branchC_18_out2_valid, branchC_18_out1_valid}), .ready_out_bus({branchC_18_out2_ready, branchC_18_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_4
		(.clk(source_4_clk), .rst(source_4_rst),
		.data_out_bus({source_4_out1_data}), .valid_out_bus({source_4_out1_valid}), .ready_out_bus({source_4_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_5
		(.clk(source_5_clk), .rst(source_5_rst),
		.data_out_bus({source_5_out1_data}), .valid_out_bus({source_5_out1_valid}), .ready_out_bus({source_5_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(6))source_node_source_6
		(.clk(source_6_clk), .rst(source_6_rst),
		.data_out_bus({source_6_out1_data}), .valid_out_bus({source_6_out1_valid}), .ready_out_bus({source_6_out1_ready}));

	ret_op #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) ret_op_ret_0
		(.clk(ret_0_clk), .rst(ret_0_rst),
		.data_in_bus({ret_0_in1_data}), .valid_in_bus({ret_0_in1_valid}), .ready_in_bus({ret_0_in1_ready}), 
		.data_out_bus({ret_0_out1_data}), .valid_out_bus({ret_0_out1_valid}), .ready_out_bus({ret_0_out1_ready}));

	end_node #(.INPUTS(1), .OUTPUTS(1), .MEMORY_INPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) end_node_end_0
		(.clk(end_0_clk), .rst(end_0_rst),
		.data_in_bus({end_0_in4_data}), .valid_in_bus({end_0_in4_valid}), .ready_in_bus({end_0_in4_ready}), .e_valid_bus({end_0_in3_valid, end_0_in2_valid, end_0_in1_valid}), .e_ready_bus({end_0_in3_ready, end_0_in2_ready, end_0_in1_ready}), 
		.data_out_bus({end_0_out1_data}), .valid_out_bus({end_0_out1_valid}), .ready_out_bus({end_0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_12
		(.clk(phiC_12_clk), .rst(phiC_12_rst),
		.data_in_bus({phiC_12_in1_data}), .valid_in_bus({phiC_12_in1_valid}), .ready_in_bus({phiC_12_in1_ready}), 
		.data_out_bus({phiC_12_out1_data}), .valid_out_bus({phiC_12_out1_valid}), .ready_out_bus({phiC_12_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6), .COND_SIZE(1)) mux_node_phi_1
		(.clk(phi_1_clk), .rst(phi_1_rst),
		.data_in_bus({{5'b0, phi_1_in1_data}, phi_1_in3_data, phi_1_in2_data}), .valid_in_bus({phi_1_in1_valid, phi_1_in3_valid, phi_1_in2_valid}), .ready_in_bus({phi_1_in1_ready, phi_1_in3_ready, phi_1_in2_ready}), 
		.data_out_bus({phi_1_out1_data}), .valid_out_bus({phi_1_out1_valid}), .ready_out_bus({phi_1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block2
		(.clk(brCst_block2_clk), .rst(brCst_block2_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block2_in1_valid}), .ready_in_bus({brCst_block2_in1_ready}), 
		.data_out_bus({brCst_block2_out1_data}), .valid_out_bus({brCst_block2_out1_valid}), .ready_out_bus({brCst_block2_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_1
		(.clk(cst_1_clk), .rst(cst_1_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_1_in1_valid}), .ready_in_bus({cst_1_in1_ready}), 
		.data_out_bus({cst_1_out1_data}), .valid_out_bus({cst_1_out1_valid}), .ready_out_bus({cst_1_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_1
		(.clk(branch_1_clk), .rst(branch_1_rst),
		.data_in_bus({{branch_1_in2_data}, branch_1_in1_data}), .valid_in_bus({branch_1_in2_valid, branch_1_in1_valid}), .ready_in_bus({branch_1_in2_ready, branch_1_in1_ready}), 
		.data_out_bus({branch_1_out2_data, branch_1_out1_data}), .valid_out_bus({branch_1_out2_valid, branch_1_out1_valid}), .ready_out_bus({branch_1_out2_ready, branch_1_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(6), .DATA_OUT_SIZE(6)) branch_node_branch_2
		(.clk(branch_2_clk), .rst(branch_2_rst),
		.data_in_bus({{5'b0, branch_2_in2_data}, branch_2_in1_data}), .valid_in_bus({branch_2_in2_valid, branch_2_in1_valid}), .ready_in_bus({branch_2_in2_ready, branch_2_in1_ready}), 
		.data_out_bus({branch_2_out2_data, branch_2_out1_data}), .valid_out_bus({branch_2_out2_valid, branch_2_out1_valid}), .ready_out_bus({branch_2_out2_ready, branch_2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_10
		(.clk(fork_10_clk), .rst(fork_10_rst),
		.data_in_bus({fork_10_in1_data}), .valid_in_bus({fork_10_in1_valid}), .ready_in_bus({fork_10_in1_ready}), 
		.data_out_bus({fork_10_out3_data, fork_10_out2_data, fork_10_out1_data}), .valid_out_bus({fork_10_out3_valid, fork_10_out2_valid, fork_10_out1_valid}), .ready_out_bus({fork_10_out3_ready, fork_10_out2_ready, fork_10_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_7
		(.clk(phiC_7_clk), .rst(phiC_7_rst),
		.data_in_bus({phiC_7_in2_data, phiC_7_in1_data}), .valid_in_bus({phiC_7_in2_valid, phiC_7_in1_valid}), .ready_in_bus({phiC_7_in2_ready, phiC_7_in1_ready}), 
		.data_out_bus({phiC_7_out2_data, phiC_7_out1_data}), .valid_out_bus({phiC_7_out2_valid, phiC_7_out1_valid}), .ready_out_bus({phiC_7_out2_ready, phiC_7_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_18
		(.clk(forkC_18_clk), .rst(forkC_18_rst),
		.data_in_bus({forkC_18_in1_data}), .valid_in_bus({forkC_18_in1_valid}), .ready_in_bus({forkC_18_in1_ready}), 
		.data_out_bus({forkC_18_out3_data, forkC_18_out2_data, forkC_18_out1_data}), .valid_out_bus({forkC_18_out3_valid, forkC_18_out2_valid, forkC_18_out1_valid}), .ready_out_bus({forkC_18_out3_ready, forkC_18_out2_ready, forkC_18_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_15
		(.clk(branchC_15_clk), .rst(branchC_15_rst),
		.data_in_bus({{branchC_15_in2_data}, branchC_15_in1_data}), .valid_in_bus({branchC_15_in2_valid, branchC_15_in1_valid}), .ready_in_bus({branchC_15_in2_ready, branchC_15_in1_ready}), 
		.data_out_bus({branchC_15_out2_data, branchC_15_out1_data}), .valid_out_bus({branchC_15_out2_valid, branchC_15_out1_valid}), .ready_out_bus({branchC_15_out2_ready, branchC_15_out1_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(12), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_in_a
		(.clk(MC_in_a_clk), .rst(MC_in_a_rst),
		.io_storeDataOut(in_a_dout0), .io_storeAddrOut(in_a_address0), .io_storeEnable(in_a_we0),
		.io_loadDataIn(in_a_din1), .io_loadAddrOut(in_a_address1), .io_loadEnable(in_a_ce1),
		.io_bbpValids({MC_in_a_in2_valid}), .io_bb_stCountArray({MC_in_a_in2_data}), .io_bbReadyToPrevs({MC_in_a_in2_ready}), .io_rdPortsPrev_ready({MC_in_a_in1_ready}), .io_rdPortsPrev_valid({MC_in_a_in1_valid}), .io_rdPortsPrev_bits({MC_in_a_in1_data}), 	
	.io_wrAddrPorts_ready({MC_in_a_in3_ready}), .io_wrAddrPorts_valid({MC_in_a_in3_valid}), .io_wrAddrPorts_bits({MC_in_a_in3_data}), 	
	.io_wrDataPorts_ready({MC_in_a_in4_ready}), .io_wrDataPorts_valid({MC_in_a_in4_valid}), .io_wrDataPorts_bits({MC_in_a_in4_data}), 	
	.io_rdPortsNext_ready({MC_in_a_out1_ready}), .io_rdPortsNext_valid({MC_in_a_out1_valid}), .io_rdPortsNext_bits({MC_in_a_out1_data}), 	
	.io_Empty_Valid({MC_in_a_out2_valid}), .io_Empty_Ready({MC_in_a_out2_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(12), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_in_b
		(.clk(MC_in_b_clk), .rst(MC_in_b_rst),
		.io_storeDataOut(in_b_dout0), .io_storeAddrOut(in_b_address0), .io_storeEnable(in_b_we0),
		.io_loadDataIn(in_b_din1), .io_loadAddrOut(in_b_address1), .io_loadEnable(in_b_ce1),
		.io_bbpValids({MC_in_b_in2_valid}), .io_bb_stCountArray({MC_in_b_in2_data}), .io_bbReadyToPrevs({MC_in_b_in2_ready}), .io_rdPortsPrev_ready({MC_in_b_in1_ready}), .io_rdPortsPrev_valid({MC_in_b_in1_valid}), .io_rdPortsPrev_bits({MC_in_b_in1_data}), 	
	.io_wrAddrPorts_ready({MC_in_b_in3_ready}), .io_wrAddrPorts_valid({MC_in_b_in3_valid}), .io_wrAddrPorts_bits({MC_in_b_in3_data}), 	
	.io_wrDataPorts_ready({MC_in_b_in4_ready}), .io_wrDataPorts_valid({MC_in_b_in4_valid}), .io_wrDataPorts_bits({MC_in_b_in4_data}), 	
	.io_rdPortsNext_ready({MC_in_b_out1_ready}), .io_rdPortsNext_valid({MC_in_b_out1_valid}), .io_rdPortsNext_bits({MC_in_b_out1_data}), 	
	.io_Empty_Valid({MC_in_b_out2_valid}), .io_Empty_Ready({MC_in_b_out2_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(12), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_out_c
		(.clk(MC_out_c_clk), .rst(MC_out_c_rst),
		.io_storeDataOut(out_c_dout0), .io_storeAddrOut(out_c_address0), .io_storeEnable(out_c_we0),
		.io_loadDataIn(out_c_din1), .io_loadAddrOut(out_c_address1), .io_loadEnable(out_c_ce1),
		.io_bbpValids({MC_out_c_in1_valid}), .io_bb_stCountArray({MC_out_c_in1_data}), .io_bbReadyToPrevs({MC_out_c_in1_ready}), .io_rdPortsPrev_ready({MC_out_c_in4_ready}), .io_rdPortsPrev_valid({MC_out_c_in4_valid}), .io_rdPortsPrev_bits({MC_out_c_in4_data}), 	
	.io_wrAddrPorts_ready({MC_out_c_in2_ready}), .io_wrAddrPorts_valid({MC_out_c_in2_valid}), .io_wrAddrPorts_bits({MC_out_c_in2_data}), 	
	.io_wrDataPorts_ready({MC_out_c_in3_ready}), .io_wrDataPorts_valid({MC_out_c_in3_valid}), .io_wrDataPorts_bits({MC_out_c_in3_data}), 	
	.io_rdPortsNext_ready({MC_out_c_out2_ready}), .io_rdPortsNext_valid({MC_out_c_out2_valid}), .io_rdPortsNext_bits({MC_out_c_out2_data}), 	
	.io_Empty_Valid({MC_out_c_out1_valid}), .io_Empty_Ready({MC_out_c_out1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_0
		(.clk(sink_0_clk), .rst(sink_0_rst),
		.data_in_bus({sink_0_in1_data}), .valid_in_bus({sink_0_in1_valid}), .ready_in_bus({sink_0_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_1
		(.clk(sink_1_clk), .rst(sink_1_rst),
		.data_in_bus({sink_1_in1_data}), .valid_in_bus({sink_1_in1_valid}), .ready_in_bus({sink_1_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_2
		(.clk(sink_2_clk), .rst(sink_2_rst),
		.data_in_bus({sink_2_in1_data}), .valid_in_bus({sink_2_in1_valid}), .ready_in_bus({sink_2_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_3
		(.clk(sink_3_clk), .rst(sink_3_rst),
		.data_in_bus({sink_3_in1_data}), .valid_in_bus({sink_3_in1_valid}), .ready_in_bus({sink_3_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_4
		(.clk(sink_4_clk), .rst(sink_4_rst),
		.data_in_bus({sink_4_in1_data}), .valid_in_bus({sink_4_in1_valid}), .ready_in_bus({sink_4_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_5
		(.clk(sink_5_clk), .rst(sink_5_rst),
		.data_in_bus({sink_5_in1_data}), .valid_in_bus({sink_5_in1_valid}), .ready_in_bus({sink_5_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_6
		(.clk(sink_6_clk), .rst(sink_6_rst),
		.data_in_bus({sink_6_in1_data}), .valid_in_bus({sink_6_in1_valid}), .ready_in_bus({sink_6_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_7
		(.clk(sink_7_clk), .rst(sink_7_rst),
		.data_in_bus({sink_7_in1_data}), .valid_in_bus({sink_7_in1_valid}), .ready_in_bus({sink_7_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_8
		(.clk(sink_8_clk), .rst(sink_8_rst),
		.data_in_bus({sink_8_in1_data}), .valid_in_bus({sink_8_in1_valid}), .ready_in_bus({sink_8_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(6))sink_node_sink_9
		(.clk(sink_9_clk), .rst(sink_9_rst),
		.data_in_bus({sink_9_in1_data}), .valid_in_bus({sink_9_in1_valid}), .ready_in_bus({sink_9_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_10
		(.clk(sink_10_clk), .rst(sink_10_rst),
		.data_in_bus({sink_10_in1_data}), .valid_in_bus({sink_10_in1_valid}), .ready_in_bus({sink_10_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_11
		(.clk(sink_11_clk), .rst(sink_11_rst),
		.data_in_bus({sink_11_in1_data}), .valid_in_bus({sink_11_in1_valid}), .ready_in_bus({sink_11_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_12
		(.clk(sink_12_clk), .rst(sink_12_rst),
		.data_in_bus({sink_12_in1_data}), .valid_in_bus({sink_12_in1_valid}), .ready_in_bus({sink_12_in1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_100
		(.clk(Buffer_100_clk), .rst(Buffer_100_rst),
		.data_in_bus({Buffer_100_in1_data}), .valid_in_bus({Buffer_100_in1_valid}), .ready_in_bus({Buffer_100_in1_ready}), 
		.data_out_bus({Buffer_100_out1_data}), .valid_out_bus({Buffer_100_out1_valid}), .ready_out_bus({Buffer_100_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_101
		(.clk(Buffer_101_clk), .rst(Buffer_101_rst),
		.data_in_bus({Buffer_101_in1_data}), .valid_in_bus({Buffer_101_in1_valid}), .ready_in_bus({Buffer_101_in1_ready}), 
		.data_out_bus({Buffer_101_out1_data}), .valid_out_bus({Buffer_101_out1_valid}), .ready_out_bus({Buffer_101_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_102
		(.clk(Buffer_102_clk), .rst(Buffer_102_rst),
		.data_in_bus({Buffer_102_in1_data}), .valid_in_bus({Buffer_102_in1_valid}), .ready_in_bus({Buffer_102_in1_ready}), 
		.data_out_bus({Buffer_102_out1_data}), .valid_out_bus({Buffer_102_out1_valid}), .ready_out_bus({Buffer_102_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_103
		(.clk(Buffer_103_clk), .rst(Buffer_103_rst),
		.data_in_bus({Buffer_103_in1_data}), .valid_in_bus({Buffer_103_in1_valid}), .ready_in_bus({Buffer_103_in1_ready}), 
		.data_out_bus({Buffer_103_out1_data}), .valid_out_bus({Buffer_103_out1_valid}), .ready_out_bus({Buffer_103_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_104
		(.clk(Buffer_104_clk), .rst(Buffer_104_rst),
		.data_in_bus({Buffer_104_in1_data}), .valid_in_bus({Buffer_104_in1_valid}), .ready_in_bus({Buffer_104_in1_ready}), 
		.data_out_bus({Buffer_104_out1_data}), .valid_out_bus({Buffer_104_out1_valid}), .ready_out_bus({Buffer_104_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_105
		(.clk(Buffer_105_clk), .rst(Buffer_105_rst),
		.data_in_bus({Buffer_105_in1_data}), .valid_in_bus({Buffer_105_in1_valid}), .ready_in_bus({Buffer_105_in1_ready}), 
		.data_out_bus({Buffer_105_out1_data}), .valid_out_bus({Buffer_105_out1_valid}), .ready_out_bus({Buffer_105_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_106
		(.clk(Buffer_106_clk), .rst(Buffer_106_rst),
		.data_in_bus({Buffer_106_in1_data}), .valid_in_bus({Buffer_106_in1_valid}), .ready_in_bus({Buffer_106_in1_ready}), 
		.data_out_bus({Buffer_106_out1_data}), .valid_out_bus({Buffer_106_out1_valid}), .ready_out_bus({Buffer_106_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_107
		(.clk(Buffer_107_clk), .rst(Buffer_107_rst),
		.data_in_bus({Buffer_107_in1_data}), .valid_in_bus({Buffer_107_in1_valid}), .ready_in_bus({Buffer_107_in1_ready}), 
		.data_out_bus({Buffer_107_out1_data}), .valid_out_bus({Buffer_107_out1_valid}), .ready_out_bus({Buffer_107_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_108
		(.clk(Buffer_108_clk), .rst(Buffer_108_rst),
		.data_in_bus({Buffer_108_in1_data}), .valid_in_bus({Buffer_108_in1_valid}), .ready_in_bus({Buffer_108_in1_ready}), 
		.data_out_bus({Buffer_108_out1_data}), .valid_out_bus({Buffer_108_out1_valid}), .ready_out_bus({Buffer_108_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_109
		(.clk(Buffer_109_clk), .rst(Buffer_109_rst),
		.data_in_bus({Buffer_109_in1_data}), .valid_in_bus({Buffer_109_in1_valid}), .ready_in_bus({Buffer_109_in1_ready}), 
		.data_out_bus({Buffer_109_out1_data}), .valid_out_bus({Buffer_109_out1_valid}), .ready_out_bus({Buffer_109_out1_ready}));

endmodule

