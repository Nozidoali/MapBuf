module kmp(
	input clk,
	input rst,

	input [0 : 0]start_in,
	input start_valid,
	output start_ready,

	output [31 : 0]end_out,
	output end_valid,
	input end_ready,

	output [31 : 0]kmpNext_address0,
	output kmpNext_ce0,
	output kmpNext_we0,
	output [31 : 0]kmpNext_dout0,
	input [31 : 0]kmpNext_din0,
	output [31 : 0]kmpNext_address1,
	output kmpNext_ce1,
	output kmpNext_we1,
	output [31 : 0]kmpNext_dout1,
	input [31 : 0]kmpNext_din1,

	output [31 : 0]pattern_address0,
	output pattern_ce0,
	output pattern_we0,
	output [31 : 0]pattern_dout0,
	input [31 : 0]pattern_din0,
	output [31 : 0]pattern_address1,
	output pattern_ce1,
	output pattern_we1,
	output [31 : 0]pattern_dout1,
	input [31 : 0]pattern_din1,

	output [9 : 0]input_address0,
	output input_ce0,
	output input_we0,
	output [31 : 0]input_dout0,
	input [31 : 0]input_din0,
	output [9 : 0]input_address1,
	output input_ce1,
	output input_we1,
	output [31 : 0]input_dout1,
	input [31 : 0]input_din1

);

	wire phi_1_clk;
	wire phi_1_rst;
	wire [0 : 0]phi_1_in1_data;
	wire phi_1_in1_ready;
	wire phi_1_in1_valid;
	wire [31 : 0]phi_1_in2_data;
	wire phi_1_in2_ready;
	wire phi_1_in2_valid;
	wire [31 : 0]phi_1_in3_data;
	wire phi_1_in3_ready;
	wire phi_1_in3_valid;
	wire [31 : 0]phi_1_out1_data;
	wire phi_1_out1_ready;
	wire phi_1_out1_valid;

	wire phi_2_clk;
	wire phi_2_rst;
	wire [0 : 0]phi_2_in1_data;
	wire phi_2_in1_ready;
	wire phi_2_in1_valid;
	wire [2 : 0]phi_2_in2_data;
	wire phi_2_in2_ready;
	wire phi_2_in2_valid;
	wire [2 : 0]phi_2_in3_data;
	wire phi_2_in3_ready;
	wire phi_2_in3_valid;
	wire [2 : 0]phi_2_out1_data;
	wire phi_2_out1_ready;
	wire phi_2_out1_valid;

	wire load_5_clk;
	wire load_5_rst;
	wire [31 : 0]load_5_in1_data;
	wire load_5_in1_ready;
	wire load_5_in1_valid;
	wire [2 : 0]load_5_in2_data;
	wire load_5_in2_ready;
	wire load_5_in2_valid;
	wire [31 : 0]load_5_out1_data;
	wire load_5_out1_ready;
	wire load_5_out1_valid;
	wire [2 : 0]load_5_out2_data;
	wire load_5_out2_ready;
	wire load_5_out2_valid;

	wire brCst_block2_clk;
	wire brCst_block2_rst;
	wire [0 : 0]brCst_block2_in1_data;
	wire brCst_block2_in1_ready;
	wire brCst_block2_in1_valid;
	wire [0 : 0]brCst_block2_out1_data;
	wire brCst_block2_out1_ready;
	wire brCst_block2_out1_valid;

	wire fork_0_clk;
	wire fork_0_rst;
	wire [2 : 0]fork_0_in1_data;
	wire fork_0_in1_ready;
	wire fork_0_in1_valid;
	wire [2 : 0]fork_0_out1_data;
	wire fork_0_out1_ready;
	wire fork_0_out1_valid;
	wire [2 : 0]fork_0_out2_data;
	wire fork_0_out2_ready;
	wire fork_0_out2_valid;

	wire branch_2_clk;
	wire branch_2_rst;
	wire [31 : 0]branch_2_in1_data;
	wire branch_2_in1_ready;
	wire branch_2_in1_valid;
	wire [0 : 0]branch_2_in2_data;
	wire branch_2_in2_ready;
	wire branch_2_in2_valid;
	wire [31 : 0]branch_2_out1_data;
	wire branch_2_out1_ready;
	wire branch_2_out1_valid;
	wire [31 : 0]branch_2_out2_data;
	wire branch_2_out2_ready;
	wire branch_2_out2_valid;

	wire branch_3_clk;
	wire branch_3_rst;
	wire [31 : 0]branch_3_in1_data;
	wire branch_3_in1_ready;
	wire branch_3_in1_valid;
	wire [0 : 0]branch_3_in2_data;
	wire branch_3_in2_ready;
	wire branch_3_in2_valid;
	wire [31 : 0]branch_3_out1_data;
	wire branch_3_out1_ready;
	wire branch_3_out1_valid;
	wire [31 : 0]branch_3_out2_data;
	wire branch_3_out2_ready;
	wire branch_3_out2_valid;

	wire branch_4_clk;
	wire branch_4_rst;
	wire [2 : 0]branch_4_in1_data;
	wire branch_4_in1_ready;
	wire branch_4_in1_valid;
	wire [0 : 0]branch_4_in2_data;
	wire branch_4_in2_ready;
	wire branch_4_in2_valid;
	wire [2 : 0]branch_4_out1_data;
	wire branch_4_out1_ready;
	wire branch_4_out1_valid;
	wire [2 : 0]branch_4_out2_data;
	wire branch_4_out2_ready;
	wire branch_4_out2_valid;

	wire fork_28_clk;
	wire fork_28_rst;
	wire [0 : 0]fork_28_in1_data;
	wire fork_28_in1_ready;
	wire fork_28_in1_valid;
	wire [0 : 0]fork_28_out1_data;
	wire fork_28_out1_ready;
	wire fork_28_out1_valid;
	wire [0 : 0]fork_28_out2_data;
	wire fork_28_out2_ready;
	wire fork_28_out2_valid;
	wire [0 : 0]fork_28_out3_data;
	wire fork_28_out3_ready;
	wire fork_28_out3_valid;
	wire [0 : 0]fork_28_out4_data;
	wire fork_28_out4_ready;
	wire fork_28_out4_valid;

	wire phiC_30_clk;
	wire phiC_30_rst;
	wire [0 : 0]phiC_30_in1_data;
	wire phiC_30_in1_ready;
	wire phiC_30_in1_valid;
	wire [0 : 0]phiC_30_in2_data;
	wire phiC_30_in2_ready;
	wire phiC_30_in2_valid;
	wire [0 : 0]phiC_30_out1_data;
	wire phiC_30_out1_ready;
	wire phiC_30_out1_valid;
	wire [0 : 0]phiC_30_out2_data;
	wire phiC_30_out2_ready;
	wire phiC_30_out2_valid;

	wire forkC_43_clk;
	wire forkC_43_rst;
	wire [0 : 0]forkC_43_in1_data;
	wire forkC_43_in1_ready;
	wire forkC_43_in1_valid;
	wire [0 : 0]forkC_43_out1_data;
	wire forkC_43_out1_ready;
	wire forkC_43_out1_valid;
	wire [0 : 0]forkC_43_out2_data;
	wire forkC_43_out2_ready;
	wire forkC_43_out2_valid;

	wire branchC_45_clk;
	wire branchC_45_rst;
	wire [0 : 0]branchC_45_in1_data;
	wire branchC_45_in1_ready;
	wire branchC_45_in1_valid;
	wire [0 : 0]branchC_45_in2_data;
	wire branchC_45_in2_ready;
	wire branchC_45_in2_valid;
	wire [0 : 0]branchC_45_out1_data;
	wire branchC_45_out1_ready;
	wire branchC_45_out1_valid;
	wire [0 : 0]branchC_45_out2_data;
	wire branchC_45_out2_ready;
	wire branchC_45_out2_valid;

	wire fork_57_clk;
	wire fork_57_rst;
	wire [0 : 0]fork_57_in1_data;
	wire fork_57_in1_ready;
	wire fork_57_in1_valid;
	wire [0 : 0]fork_57_out1_data;
	wire fork_57_out1_ready;
	wire fork_57_out1_valid;
	wire [0 : 0]fork_57_out2_data;
	wire fork_57_out2_ready;
	wire fork_57_out2_valid;

	wire phi_31_clk;
	wire phi_31_rst;
	wire [0 : 0]phi_31_in1_data;
	wire phi_31_in1_ready;
	wire phi_31_in1_valid;
	wire [31 : 0]phi_31_in2_data;
	wire phi_31_in2_ready;
	wire phi_31_in2_valid;
	wire [31 : 0]phi_31_in3_data;
	wire phi_31_in3_ready;
	wire phi_31_in3_valid;
	wire [31 : 0]phi_31_out1_data;
	wire phi_31_out1_ready;
	wire phi_31_out1_valid;

	wire phi_32_clk;
	wire phi_32_rst;
	wire [0 : 0]phi_32_in1_data;
	wire phi_32_in1_ready;
	wire phi_32_in1_valid;
	wire [31 : 0]phi_32_in2_data;
	wire phi_32_in2_ready;
	wire phi_32_in2_valid;
	wire [31 : 0]phi_32_in3_data;
	wire phi_32_in3_ready;
	wire phi_32_in3_valid;
	wire [31 : 0]phi_32_out1_data;
	wire phi_32_out1_ready;
	wire phi_32_out1_valid;

	wire phi_33_clk;
	wire phi_33_rst;
	wire [0 : 0]phi_33_in1_data;
	wire phi_33_in1_ready;
	wire phi_33_in1_valid;
	wire [9 : 0]phi_33_in2_data;
	wire phi_33_in2_ready;
	wire phi_33_in2_valid;
	wire [9 : 0]phi_33_in3_data;
	wire phi_33_in3_ready;
	wire phi_33_in3_valid;
	wire [9 : 0]phi_33_out1_data;
	wire phi_33_out1_ready;
	wire phi_33_out1_valid;

	wire load_36_clk;
	wire load_36_rst;
	wire [31 : 0]load_36_in1_data;
	wire load_36_in1_ready;
	wire load_36_in1_valid;
	wire [9 : 0]load_36_in2_data;
	wire load_36_in2_ready;
	wire load_36_in2_valid;
	wire [31 : 0]load_36_out1_data;
	wire load_36_out1_ready;
	wire load_36_out1_valid;
	wire [9 : 0]load_36_out2_data;
	wire load_36_out2_ready;
	wire load_36_out2_valid;

	wire brCst_block8_clk;
	wire brCst_block8_rst;
	wire [0 : 0]brCst_block8_in1_data;
	wire brCst_block8_in1_ready;
	wire brCst_block8_in1_valid;
	wire [0 : 0]brCst_block8_out1_data;
	wire brCst_block8_out1_ready;
	wire brCst_block8_out1_valid;

	wire fork_4_clk;
	wire fork_4_rst;
	wire [9 : 0]fork_4_in1_data;
	wire fork_4_in1_ready;
	wire fork_4_in1_valid;
	wire [9 : 0]fork_4_out1_data;
	wire fork_4_out1_ready;
	wire fork_4_out1_valid;
	wire [9 : 0]fork_4_out2_data;
	wire fork_4_out2_ready;
	wire fork_4_out2_valid;

	wire branch_19_clk;
	wire branch_19_rst;
	wire [31 : 0]branch_19_in1_data;
	wire branch_19_in1_ready;
	wire branch_19_in1_valid;
	wire [0 : 0]branch_19_in2_data;
	wire branch_19_in2_ready;
	wire branch_19_in2_valid;
	wire [31 : 0]branch_19_out1_data;
	wire branch_19_out1_ready;
	wire branch_19_out1_valid;
	wire [31 : 0]branch_19_out2_data;
	wire branch_19_out2_ready;
	wire branch_19_out2_valid;

	wire branch_20_clk;
	wire branch_20_rst;
	wire [31 : 0]branch_20_in1_data;
	wire branch_20_in1_ready;
	wire branch_20_in1_valid;
	wire [0 : 0]branch_20_in2_data;
	wire branch_20_in2_ready;
	wire branch_20_in2_valid;
	wire [31 : 0]branch_20_out1_data;
	wire branch_20_out1_ready;
	wire branch_20_out1_valid;
	wire [31 : 0]branch_20_out2_data;
	wire branch_20_out2_ready;
	wire branch_20_out2_valid;

	wire branch_21_clk;
	wire branch_21_rst;
	wire [31 : 0]branch_21_in1_data;
	wire branch_21_in1_ready;
	wire branch_21_in1_valid;
	wire [0 : 0]branch_21_in2_data;
	wire branch_21_in2_ready;
	wire branch_21_in2_valid;
	wire [31 : 0]branch_21_out1_data;
	wire branch_21_out1_ready;
	wire branch_21_out1_valid;
	wire [31 : 0]branch_21_out2_data;
	wire branch_21_out2_ready;
	wire branch_21_out2_valid;

	wire branch_22_clk;
	wire branch_22_rst;
	wire [9 : 0]branch_22_in1_data;
	wire branch_22_in1_ready;
	wire branch_22_in1_valid;
	wire [0 : 0]branch_22_in2_data;
	wire branch_22_in2_ready;
	wire branch_22_in2_valid;
	wire [9 : 0]branch_22_out1_data;
	wire branch_22_out1_ready;
	wire branch_22_out1_valid;
	wire [9 : 0]branch_22_out2_data;
	wire branch_22_out2_ready;
	wire branch_22_out2_valid;

	wire fork_34_clk;
	wire fork_34_rst;
	wire [0 : 0]fork_34_in1_data;
	wire fork_34_in1_ready;
	wire fork_34_in1_valid;
	wire [0 : 0]fork_34_out1_data;
	wire fork_34_out1_ready;
	wire fork_34_out1_valid;
	wire [0 : 0]fork_34_out2_data;
	wire fork_34_out2_ready;
	wire fork_34_out2_valid;
	wire [0 : 0]fork_34_out3_data;
	wire fork_34_out3_ready;
	wire fork_34_out3_valid;
	wire [0 : 0]fork_34_out4_data;
	wire fork_34_out4_ready;
	wire fork_34_out4_valid;
	wire [0 : 0]fork_34_out5_data;
	wire fork_34_out5_ready;
	wire fork_34_out5_valid;

	wire phiC_36_clk;
	wire phiC_36_rst;
	wire [0 : 0]phiC_36_in1_data;
	wire phiC_36_in1_ready;
	wire phiC_36_in1_valid;
	wire [0 : 0]phiC_36_in2_data;
	wire phiC_36_in2_ready;
	wire phiC_36_in2_valid;
	wire [0 : 0]phiC_36_out1_data;
	wire phiC_36_out1_ready;
	wire phiC_36_out1_valid;
	wire [0 : 0]phiC_36_out2_data;
	wire phiC_36_out2_ready;
	wire phiC_36_out2_valid;

	wire forkC_49_clk;
	wire forkC_49_rst;
	wire [0 : 0]forkC_49_in1_data;
	wire forkC_49_in1_ready;
	wire forkC_49_in1_valid;
	wire [0 : 0]forkC_49_out1_data;
	wire forkC_49_out1_ready;
	wire forkC_49_out1_valid;
	wire [0 : 0]forkC_49_out2_data;
	wire forkC_49_out2_ready;
	wire forkC_49_out2_valid;

	wire branchC_51_clk;
	wire branchC_51_rst;
	wire [0 : 0]branchC_51_in1_data;
	wire branchC_51_in1_ready;
	wire branchC_51_in1_valid;
	wire [0 : 0]branchC_51_in2_data;
	wire branchC_51_in2_ready;
	wire branchC_51_in2_valid;
	wire [0 : 0]branchC_51_out1_data;
	wire branchC_51_out1_ready;
	wire branchC_51_out1_valid;
	wire [0 : 0]branchC_51_out2_data;
	wire branchC_51_out2_ready;
	wire branchC_51_out2_valid;

	wire fork_59_clk;
	wire fork_59_rst;
	wire [0 : 0]fork_59_in1_data;
	wire fork_59_in1_ready;
	wire fork_59_in1_valid;
	wire [0 : 0]fork_59_out1_data;
	wire fork_59_out1_ready;
	wire fork_59_out1_valid;
	wire [0 : 0]fork_59_out2_data;
	wire fork_59_out2_ready;
	wire fork_59_out2_valid;
	wire [0 : 0]fork_59_out3_data;
	wire fork_59_out3_ready;
	wire fork_59_out3_valid;

	wire load_48_clk;
	wire load_48_rst;
	wire [31 : 0]load_48_in1_data;
	wire load_48_in1_ready;
	wire load_48_in1_valid;
	wire [31 : 0]load_48_in2_data;
	wire load_48_in2_ready;
	wire load_48_in2_valid;
	wire [31 : 0]load_48_out1_data;
	wire load_48_out1_ready;
	wire load_48_out1_valid;
	wire [31 : 0]load_48_out2_data;
	wire load_48_out2_ready;
	wire load_48_out2_valid;

	wire brCst_block11_clk;
	wire brCst_block11_rst;
	wire [0 : 0]brCst_block11_in1_data;
	wire brCst_block11_in1_ready;
	wire brCst_block11_in1_valid;
	wire [0 : 0]brCst_block11_out1_data;
	wire brCst_block11_out1_ready;
	wire brCst_block11_out1_valid;

	wire phi_n17_clk;
	wire phi_n17_rst;
	wire [31 : 0]phi_n17_in1_data;
	wire phi_n17_in1_ready;
	wire phi_n17_in1_valid;
	wire [31 : 0]phi_n17_out1_data;
	wire phi_n17_out1_ready;
	wire phi_n17_out1_valid;

	wire phi_n18_clk;
	wire phi_n18_rst;
	wire [31 : 0]phi_n18_in1_data;
	wire phi_n18_in1_ready;
	wire phi_n18_in1_valid;
	wire [31 : 0]phi_n18_out1_data;
	wire phi_n18_out1_ready;
	wire phi_n18_out1_valid;

	wire phi_n19_clk;
	wire phi_n19_rst;
	wire [31 : 0]phi_n19_in1_data;
	wire phi_n19_in1_ready;
	wire phi_n19_in1_valid;
	wire [31 : 0]phi_n19_out1_data;
	wire phi_n19_out1_ready;
	wire phi_n19_out1_valid;

	wire phi_n20_clk;
	wire phi_n20_rst;
	wire [9 : 0]phi_n20_in1_data;
	wire phi_n20_in1_ready;
	wire phi_n20_in1_valid;
	wire [9 : 0]phi_n20_out1_data;
	wire phi_n20_out1_ready;
	wire phi_n20_out1_valid;

	wire branch_31_clk;
	wire branch_31_rst;
	wire [31 : 0]branch_31_in1_data;
	wire branch_31_in1_ready;
	wire branch_31_in1_valid;
	wire [0 : 0]branch_31_in2_data;
	wire branch_31_in2_ready;
	wire branch_31_in2_valid;
	wire [31 : 0]branch_31_out1_data;
	wire branch_31_out1_ready;
	wire branch_31_out1_valid;
	wire [31 : 0]branch_31_out2_data;
	wire branch_31_out2_ready;
	wire branch_31_out2_valid;

	wire branch_32_clk;
	wire branch_32_rst;
	wire [31 : 0]branch_32_in1_data;
	wire branch_32_in1_ready;
	wire branch_32_in1_valid;
	wire [0 : 0]branch_32_in2_data;
	wire branch_32_in2_ready;
	wire branch_32_in2_valid;
	wire [31 : 0]branch_32_out1_data;
	wire branch_32_out1_ready;
	wire branch_32_out1_valid;
	wire [31 : 0]branch_32_out2_data;
	wire branch_32_out2_ready;
	wire branch_32_out2_valid;

	wire branch_33_clk;
	wire branch_33_rst;
	wire [31 : 0]branch_33_in1_data;
	wire branch_33_in1_ready;
	wire branch_33_in1_valid;
	wire [0 : 0]branch_33_in2_data;
	wire branch_33_in2_ready;
	wire branch_33_in2_valid;
	wire [31 : 0]branch_33_out1_data;
	wire branch_33_out1_ready;
	wire branch_33_out1_valid;
	wire [31 : 0]branch_33_out2_data;
	wire branch_33_out2_ready;
	wire branch_33_out2_valid;

	wire branch_34_clk;
	wire branch_34_rst;
	wire [9 : 0]branch_34_in1_data;
	wire branch_34_in1_ready;
	wire branch_34_in1_valid;
	wire [0 : 0]branch_34_in2_data;
	wire branch_34_in2_ready;
	wire branch_34_in2_valid;
	wire [9 : 0]branch_34_out1_data;
	wire branch_34_out1_ready;
	wire branch_34_out1_valid;
	wire [9 : 0]branch_34_out2_data;
	wire branch_34_out2_ready;
	wire branch_34_out2_valid;

	wire fork_37_clk;
	wire fork_37_rst;
	wire [0 : 0]fork_37_in1_data;
	wire fork_37_in1_ready;
	wire fork_37_in1_valid;
	wire [0 : 0]fork_37_out1_data;
	wire fork_37_out1_ready;
	wire fork_37_out1_valid;
	wire [0 : 0]fork_37_out2_data;
	wire fork_37_out2_ready;
	wire fork_37_out2_valid;
	wire [0 : 0]fork_37_out3_data;
	wire fork_37_out3_ready;
	wire fork_37_out3_valid;
	wire [0 : 0]fork_37_out4_data;
	wire fork_37_out4_ready;
	wire fork_37_out4_valid;
	wire [0 : 0]fork_37_out5_data;
	wire fork_37_out5_ready;
	wire fork_37_out5_valid;

	wire phiC_39_clk;
	wire phiC_39_rst;
	wire [0 : 0]phiC_39_in1_data;
	wire phiC_39_in1_ready;
	wire phiC_39_in1_valid;
	wire [0 : 0]phiC_39_out1_data;
	wire phiC_39_out1_ready;
	wire phiC_39_out1_valid;

	wire forkC_52_clk;
	wire forkC_52_rst;
	wire [0 : 0]forkC_52_in1_data;
	wire forkC_52_in1_ready;
	wire forkC_52_in1_valid;
	wire [0 : 0]forkC_52_out1_data;
	wire forkC_52_out1_ready;
	wire forkC_52_out1_valid;
	wire [0 : 0]forkC_52_out2_data;
	wire forkC_52_out2_ready;
	wire forkC_52_out2_valid;

	wire branchC_54_clk;
	wire branchC_54_rst;
	wire [0 : 0]branchC_54_in1_data;
	wire branchC_54_in1_ready;
	wire branchC_54_in1_valid;
	wire [0 : 0]branchC_54_in2_data;
	wire branchC_54_in2_ready;
	wire branchC_54_in2_valid;
	wire [0 : 0]branchC_54_out1_data;
	wire branchC_54_out1_ready;
	wire branchC_54_out1_valid;
	wire [0 : 0]branchC_54_out2_data;
	wire branchC_54_out2_ready;
	wire branchC_54_out2_valid;

	wire load_52_clk;
	wire load_52_rst;
	wire [31 : 0]load_52_in1_data;
	wire load_52_in1_ready;
	wire load_52_in1_valid;
	wire [31 : 0]load_52_in2_data;
	wire load_52_in2_ready;
	wire load_52_in2_valid;
	wire [31 : 0]load_52_out1_data;
	wire load_52_out1_ready;
	wire load_52_out1_valid;
	wire [31 : 0]load_52_out2_data;
	wire load_52_out2_ready;
	wire load_52_out2_valid;

	wire icmp_53_clk;
	wire icmp_53_rst;
	wire [31 : 0]icmp_53_in1_data;
	wire icmp_53_in1_ready;
	wire icmp_53_in1_valid;
	wire [31 : 0]icmp_53_in2_data;
	wire icmp_53_in2_ready;
	wire icmp_53_in2_valid;
	wire [0 : 0]icmp_53_out1_data;
	wire icmp_53_out1_ready;
	wire icmp_53_out1_valid;

	wire zext_54_clk;
	wire zext_54_rst;
	wire [0 : 0]zext_54_in1_data;
	wire zext_54_in1_ready;
	wire zext_54_in1_valid;
	wire [0 : 0]zext_54_out1_data;
	wire zext_54_out1_ready;
	wire zext_54_out1_valid;

	wire add_55_clk;
	wire add_55_rst;
	wire [31 : 0]add_55_in1_data;
	wire add_55_in1_ready;
	wire add_55_in1_valid;
	wire [31 : 0]add_55_in2_data;
	wire add_55_in2_ready;
	wire add_55_in2_valid;
	wire [31 : 0]add_55_out1_data;
	wire add_55_out1_ready;
	wire add_55_out1_valid;

	wire cst_10_clk;
	wire cst_10_rst;
	wire [1 : 0]cst_10_in1_data;
	wire cst_10_in1_ready;
	wire cst_10_in1_valid;
	wire [1 : 0]cst_10_out1_data;
	wire cst_10_out1_ready;
	wire cst_10_out1_valid;

	wire icmp_56_clk;
	wire icmp_56_rst;
	wire [31 : 0]icmp_56_in1_data;
	wire icmp_56_in1_ready;
	wire icmp_56_in1_valid;
	wire [31 : 0]icmp_56_in2_data;
	wire icmp_56_in2_ready;
	wire icmp_56_in2_valid;
	wire [0 : 0]icmp_56_out1_data;
	wire icmp_56_out1_ready;
	wire icmp_56_out1_valid;

	wire phi_n25_clk;
	wire phi_n25_rst;
	wire [31 : 0]phi_n25_in1_data;
	wire phi_n25_in1_ready;
	wire phi_n25_in1_valid;
	wire [31 : 0]phi_n25_in2_data;
	wire phi_n25_in2_ready;
	wire phi_n25_in2_valid;
	wire [31 : 0]phi_n25_out1_data;
	wire phi_n25_out1_ready;
	wire phi_n25_out1_valid;

	wire phi_n26_clk;
	wire phi_n26_rst;
	wire [31 : 0]phi_n26_in1_data;
	wire phi_n26_in1_ready;
	wire phi_n26_in1_valid;
	wire [31 : 0]phi_n26_in2_data;
	wire phi_n26_in2_ready;
	wire phi_n26_in2_valid;
	wire [31 : 0]phi_n26_out1_data;
	wire phi_n26_out1_ready;
	wire phi_n26_out1_valid;

	wire phi_n27_clk;
	wire phi_n27_rst;
	wire [31 : 0]phi_n27_in1_data;
	wire phi_n27_in1_ready;
	wire phi_n27_in1_valid;
	wire [31 : 0]phi_n27_in2_data;
	wire phi_n27_in2_ready;
	wire phi_n27_in2_valid;
	wire [31 : 0]phi_n27_out1_data;
	wire phi_n27_out1_ready;
	wire phi_n27_out1_valid;

	wire phi_n28_clk;
	wire phi_n28_rst;
	wire [9 : 0]phi_n28_in1_data;
	wire phi_n28_in1_ready;
	wire phi_n28_in1_valid;
	wire [9 : 0]phi_n28_in2_data;
	wire phi_n28_in2_ready;
	wire phi_n28_in2_valid;
	wire [9 : 0]phi_n28_out1_data;
	wire phi_n28_out1_ready;
	wire phi_n28_out1_valid;

	wire fork_6_clk;
	wire fork_6_rst;
	wire [31 : 0]fork_6_in1_data;
	wire fork_6_in1_ready;
	wire fork_6_in1_valid;
	wire [31 : 0]fork_6_out1_data;
	wire fork_6_out1_ready;
	wire fork_6_out1_valid;
	wire [31 : 0]fork_6_out2_data;
	wire fork_6_out2_ready;
	wire fork_6_out2_valid;

	wire fork_24_clk;
	wire fork_24_rst;
	wire [31 : 0]fork_24_in1_data;
	wire fork_24_in1_ready;
	wire fork_24_in1_valid;
	wire [31 : 0]fork_24_out1_data;
	wire fork_24_out1_ready;
	wire fork_24_out1_valid;
	wire [31 : 0]fork_24_out2_data;
	wire fork_24_out2_ready;
	wire fork_24_out2_valid;

	wire branch_35_clk;
	wire branch_35_rst;
	wire [31 : 0]branch_35_in1_data;
	wire branch_35_in1_ready;
	wire branch_35_in1_valid;
	wire [0 : 0]branch_35_in2_data;
	wire branch_35_in2_ready;
	wire branch_35_in2_valid;
	wire [31 : 0]branch_35_out1_data;
	wire branch_35_out1_ready;
	wire branch_35_out1_valid;
	wire [31 : 0]branch_35_out2_data;
	wire branch_35_out2_ready;
	wire branch_35_out2_valid;

	wire branch_36_clk;
	wire branch_36_rst;
	wire [31 : 0]branch_36_in1_data;
	wire branch_36_in1_ready;
	wire branch_36_in1_valid;
	wire [0 : 0]branch_36_in2_data;
	wire branch_36_in2_ready;
	wire branch_36_in2_valid;
	wire [31 : 0]branch_36_out1_data;
	wire branch_36_out1_ready;
	wire branch_36_out1_valid;
	wire [31 : 0]branch_36_out2_data;
	wire branch_36_out2_ready;
	wire branch_36_out2_valid;

	wire branch_37_clk;
	wire branch_37_rst;
	wire [9 : 0]branch_37_in1_data;
	wire branch_37_in1_ready;
	wire branch_37_in1_valid;
	wire [0 : 0]branch_37_in2_data;
	wire branch_37_in2_ready;
	wire branch_37_in2_valid;
	wire [9 : 0]branch_37_out1_data;
	wire branch_37_out1_ready;
	wire branch_37_out1_valid;
	wire [9 : 0]branch_37_out2_data;
	wire branch_37_out2_ready;
	wire branch_37_out2_valid;

	wire fork_38_clk;
	wire fork_38_rst;
	wire [0 : 0]fork_38_in1_data;
	wire fork_38_in1_ready;
	wire fork_38_in1_valid;
	wire [0 : 0]fork_38_out1_data;
	wire fork_38_out1_ready;
	wire fork_38_out1_valid;
	wire [0 : 0]fork_38_out2_data;
	wire fork_38_out2_ready;
	wire fork_38_out2_valid;
	wire [0 : 0]fork_38_out3_data;
	wire fork_38_out3_ready;
	wire fork_38_out3_valid;
	wire [0 : 0]fork_38_out4_data;
	wire fork_38_out4_ready;
	wire fork_38_out4_valid;

	wire phiC_40_clk;
	wire phiC_40_rst;
	wire [0 : 0]phiC_40_in1_data;
	wire phiC_40_in1_ready;
	wire phiC_40_in1_valid;
	wire [0 : 0]phiC_40_in2_data;
	wire phiC_40_in2_ready;
	wire phiC_40_in2_valid;
	wire [0 : 0]phiC_40_out1_data;
	wire phiC_40_out1_ready;
	wire phiC_40_out1_valid;

	wire branchC_55_clk;
	wire branchC_55_rst;
	wire [0 : 0]branchC_55_in1_data;
	wire branchC_55_in1_ready;
	wire branchC_55_in1_valid;
	wire [0 : 0]branchC_55_in2_data;
	wire branchC_55_in2_ready;
	wire branchC_55_in2_valid;
	wire [0 : 0]branchC_55_out1_data;
	wire branchC_55_out1_ready;
	wire branchC_55_out1_valid;
	wire [0 : 0]branchC_55_out2_data;
	wire branchC_55_out2_ready;
	wire branchC_55_out2_valid;

	wire source_4_clk;
	wire source_4_rst;
	wire [1 : 0]source_4_out1_data;
	wire source_4_out1_ready;
	wire source_4_out1_valid;

	wire cst_0_clk;
	wire cst_0_rst;
	wire [0 : 0]cst_0_in1_data;
	wire cst_0_in1_ready;
	wire cst_0_in1_valid;
	wire [0 : 0]cst_0_out1_data;
	wire cst_0_out1_ready;
	wire cst_0_out1_valid;

	wire store_0_clk;
	wire store_0_rst;
	wire [0 : 0]store_0_in1_data;
	wire store_0_in1_ready;
	wire store_0_in1_valid;
	wire [0 : 0]store_0_in2_data;
	wire store_0_in2_ready;
	wire store_0_in2_valid;
	wire [0 : 0]store_0_out1_data;
	wire store_0_out1_ready;
	wire store_0_out1_valid;
	wire [0 : 0]store_0_out2_data;
	wire store_0_out2_ready;
	wire store_0_out2_valid;

	wire brCst_block1_clk;
	wire brCst_block1_rst;
	wire [0 : 0]brCst_block1_in1_data;
	wire brCst_block1_in1_ready;
	wire brCst_block1_in1_valid;
	wire [0 : 0]brCst_block1_out1_data;
	wire brCst_block1_out1_ready;
	wire brCst_block1_out1_valid;

	wire cst_1_clk;
	wire cst_1_rst;
	wire [0 : 0]cst_1_in1_data;
	wire cst_1_in1_ready;
	wire cst_1_in1_valid;
	wire [0 : 0]cst_1_out1_data;
	wire cst_1_out1_ready;
	wire cst_1_out1_valid;

	wire cst_2_clk;
	wire cst_2_rst;
	wire [0 : 0]cst_2_in1_data;
	wire cst_2_in1_ready;
	wire cst_2_in1_valid;
	wire [0 : 0]cst_2_out1_data;
	wire cst_2_out1_ready;
	wire cst_2_out1_valid;

	wire cst_15_clk;
	wire cst_15_rst;
	wire [0 : 0]cst_15_in1_data;
	wire cst_15_in1_ready;
	wire cst_15_in1_valid;
	wire [0 : 0]cst_15_out1_data;
	wire cst_15_out1_ready;
	wire cst_15_out1_valid;

	wire branch_0_clk;
	wire branch_0_rst;
	wire [0 : 0]branch_0_in1_data;
	wire branch_0_in1_ready;
	wire branch_0_in1_valid;
	wire [0 : 0]branch_0_in2_data;
	wire branch_0_in2_ready;
	wire branch_0_in2_valid;
	wire [0 : 0]branch_0_out1_data;
	wire branch_0_out1_ready;
	wire branch_0_out1_valid;
	wire [0 : 0]branch_0_out2_data;
	wire branch_0_out2_ready;
	wire branch_0_out2_valid;

	wire branch_1_clk;
	wire branch_1_rst;
	wire [0 : 0]branch_1_in1_data;
	wire branch_1_in1_ready;
	wire branch_1_in1_valid;
	wire [0 : 0]branch_1_in2_data;
	wire branch_1_in2_ready;
	wire branch_1_in2_valid;
	wire [0 : 0]branch_1_out1_data;
	wire branch_1_out1_ready;
	wire branch_1_out1_valid;
	wire [0 : 0]branch_1_out2_data;
	wire branch_1_out2_ready;
	wire branch_1_out2_valid;

	wire fork_27_clk;
	wire fork_27_rst;
	wire [0 : 0]fork_27_in1_data;
	wire fork_27_in1_ready;
	wire fork_27_in1_valid;
	wire [0 : 0]fork_27_out1_data;
	wire fork_27_out1_ready;
	wire fork_27_out1_valid;
	wire [0 : 0]fork_27_out2_data;
	wire fork_27_out2_ready;
	wire fork_27_out2_valid;
	wire [0 : 0]fork_27_out3_data;
	wire fork_27_out3_ready;
	wire fork_27_out3_valid;

	wire cst_16_clk;
	wire cst_16_rst;
	wire [0 : 0]cst_16_in1_data;
	wire cst_16_in1_ready;
	wire cst_16_in1_valid;
	wire [0 : 0]cst_16_out1_data;
	wire cst_16_out1_ready;
	wire cst_16_out1_valid;

	wire start_0_clk;
	wire start_0_rst;
	wire [0 : 0]start_0_in1_data;
	wire start_0_in1_ready;
	wire start_0_in1_valid;
	wire [0 : 0]start_0_out1_data;
	wire start_0_out1_ready;
	wire start_0_out1_valid;

	wire forkC_42_clk;
	wire forkC_42_rst;
	wire [0 : 0]forkC_42_in1_data;
	wire forkC_42_in1_ready;
	wire forkC_42_in1_valid;
	wire [0 : 0]forkC_42_out1_data;
	wire forkC_42_out1_ready;
	wire forkC_42_out1_valid;
	wire [0 : 0]forkC_42_out2_data;
	wire forkC_42_out2_ready;
	wire forkC_42_out2_valid;
	wire [0 : 0]forkC_42_out3_data;
	wire forkC_42_out3_ready;
	wire forkC_42_out3_valid;
	wire [0 : 0]forkC_42_out4_data;
	wire forkC_42_out4_ready;
	wire forkC_42_out4_valid;
	wire [0 : 0]forkC_42_out5_data;
	wire forkC_42_out5_ready;
	wire forkC_42_out5_valid;
	wire [0 : 0]forkC_42_out6_data;
	wire forkC_42_out6_ready;
	wire forkC_42_out6_valid;
	wire [0 : 0]forkC_42_out7_data;
	wire forkC_42_out7_ready;
	wire forkC_42_out7_valid;

	wire branchC_44_clk;
	wire branchC_44_rst;
	wire [0 : 0]branchC_44_in1_data;
	wire branchC_44_in1_ready;
	wire branchC_44_in1_valid;
	wire [0 : 0]branchC_44_in2_data;
	wire branchC_44_in2_ready;
	wire branchC_44_in2_valid;
	wire [0 : 0]branchC_44_out1_data;
	wire branchC_44_out1_ready;
	wire branchC_44_out1_valid;
	wire [0 : 0]branchC_44_out2_data;
	wire branchC_44_out2_ready;
	wire branchC_44_out2_valid;

	wire brCst_block7_clk;
	wire brCst_block7_rst;
	wire [0 : 0]brCst_block7_in1_data;
	wire brCst_block7_in1_ready;
	wire brCst_block7_in1_valid;
	wire [0 : 0]brCst_block7_out1_data;
	wire brCst_block7_out1_ready;
	wire brCst_block7_out1_valid;

	wire cst_6_clk;
	wire cst_6_rst;
	wire [0 : 0]cst_6_in1_data;
	wire cst_6_in1_ready;
	wire cst_6_in1_valid;
	wire [0 : 0]cst_6_out1_data;
	wire cst_6_out1_ready;
	wire cst_6_out1_valid;

	wire cst_7_clk;
	wire cst_7_rst;
	wire [0 : 0]cst_7_in1_data;
	wire cst_7_in1_ready;
	wire cst_7_in1_valid;
	wire [0 : 0]cst_7_out1_data;
	wire cst_7_out1_ready;
	wire cst_7_out1_valid;

	wire cst_8_clk;
	wire cst_8_rst;
	wire [0 : 0]cst_8_in1_data;
	wire cst_8_in1_ready;
	wire cst_8_in1_valid;
	wire [0 : 0]cst_8_out1_data;
	wire cst_8_out1_ready;
	wire cst_8_out1_valid;

	wire branch_16_clk;
	wire branch_16_rst;
	wire [0 : 0]branch_16_in1_data;
	wire branch_16_in1_ready;
	wire branch_16_in1_valid;
	wire [0 : 0]branch_16_in2_data;
	wire branch_16_in2_ready;
	wire branch_16_in2_valid;
	wire [0 : 0]branch_16_out1_data;
	wire branch_16_out1_ready;
	wire branch_16_out1_valid;
	wire [0 : 0]branch_16_out2_data;
	wire branch_16_out2_ready;
	wire branch_16_out2_valid;

	wire branch_17_clk;
	wire branch_17_rst;
	wire [0 : 0]branch_17_in1_data;
	wire branch_17_in1_ready;
	wire branch_17_in1_valid;
	wire [0 : 0]branch_17_in2_data;
	wire branch_17_in2_ready;
	wire branch_17_in2_valid;
	wire [0 : 0]branch_17_out1_data;
	wire branch_17_out1_ready;
	wire branch_17_out1_valid;
	wire [0 : 0]branch_17_out2_data;
	wire branch_17_out2_ready;
	wire branch_17_out2_valid;

	wire branch_18_clk;
	wire branch_18_rst;
	wire [0 : 0]branch_18_in1_data;
	wire branch_18_in1_ready;
	wire branch_18_in1_valid;
	wire [0 : 0]branch_18_in2_data;
	wire branch_18_in2_ready;
	wire branch_18_in2_valid;
	wire [0 : 0]branch_18_out1_data;
	wire branch_18_out1_ready;
	wire branch_18_out1_valid;
	wire [0 : 0]branch_18_out2_data;
	wire branch_18_out2_ready;
	wire branch_18_out2_valid;

	wire fork_33_clk;
	wire fork_33_rst;
	wire [0 : 0]fork_33_in1_data;
	wire fork_33_in1_ready;
	wire fork_33_in1_valid;
	wire [0 : 0]fork_33_out1_data;
	wire fork_33_out1_ready;
	wire fork_33_out1_valid;
	wire [0 : 0]fork_33_out2_data;
	wire fork_33_out2_ready;
	wire fork_33_out2_valid;
	wire [0 : 0]fork_33_out3_data;
	wire fork_33_out3_ready;
	wire fork_33_out3_valid;
	wire [0 : 0]fork_33_out4_data;
	wire fork_33_out4_ready;
	wire fork_33_out4_valid;

	wire phiC_35_clk;
	wire phiC_35_rst;
	wire [0 : 0]phiC_35_in1_data;
	wire phiC_35_in1_ready;
	wire phiC_35_in1_valid;
	wire [0 : 0]phiC_35_out1_data;
	wire phiC_35_out1_ready;
	wire phiC_35_out1_valid;

	wire forkC_48_clk;
	wire forkC_48_rst;
	wire [0 : 0]forkC_48_in1_data;
	wire forkC_48_in1_ready;
	wire forkC_48_in1_valid;
	wire [0 : 0]forkC_48_out1_data;
	wire forkC_48_out1_ready;
	wire forkC_48_out1_valid;
	wire [0 : 0]forkC_48_out2_data;
	wire forkC_48_out2_ready;
	wire forkC_48_out2_valid;
	wire [0 : 0]forkC_48_out3_data;
	wire forkC_48_out3_ready;
	wire forkC_48_out3_valid;
	wire [0 : 0]forkC_48_out4_data;
	wire forkC_48_out4_ready;
	wire forkC_48_out4_valid;
	wire [0 : 0]forkC_48_out5_data;
	wire forkC_48_out5_ready;
	wire forkC_48_out5_valid;

	wire branchC_50_clk;
	wire branchC_50_rst;
	wire [0 : 0]branchC_50_in1_data;
	wire branchC_50_in1_ready;
	wire branchC_50_in1_valid;
	wire [0 : 0]branchC_50_in2_data;
	wire branchC_50_in2_ready;
	wire branchC_50_in2_valid;
	wire [0 : 0]branchC_50_out1_data;
	wire branchC_50_out1_ready;
	wire branchC_50_out1_valid;
	wire [0 : 0]branchC_50_out2_data;
	wire branchC_50_out2_ready;
	wire branchC_50_out2_valid;

	wire ret_0_clk;
	wire ret_0_rst;
	wire [31 : 0]ret_0_in1_data;
	wire ret_0_in1_ready;
	wire ret_0_in1_valid;
	wire [31 : 0]ret_0_out1_data;
	wire ret_0_out1_ready;
	wire ret_0_out1_valid;

	wire phi_n29_clk;
	wire phi_n29_rst;
	wire [31 : 0]phi_n29_in1_data;
	wire phi_n29_in1_ready;
	wire phi_n29_in1_valid;
	wire [31 : 0]phi_n29_out1_data;
	wire phi_n29_out1_ready;
	wire phi_n29_out1_valid;

	wire end_0_clk;
	wire end_0_rst;
	wire [0 : 0]end_0_in1_data;
	wire end_0_in1_ready;
	wire end_0_in1_valid;
	wire [0 : 0]end_0_in2_data;
	wire end_0_in2_ready;
	wire end_0_in2_valid;
	wire [0 : 0]end_0_in3_data;
	wire end_0_in3_ready;
	wire end_0_in3_valid;
	wire [31 : 0]end_0_in4_data;
	wire end_0_in4_ready;
	wire end_0_in4_valid;
	wire [31 : 0]end_0_out1_data;
	wire end_0_out1_ready;
	wire end_0_out1_valid;

	wire phiC_43_clk;
	wire phiC_43_rst;
	wire [0 : 0]phiC_43_in1_data;
	wire phiC_43_in1_ready;
	wire phiC_43_in1_valid;
	wire [0 : 0]phiC_43_out1_data;
	wire phiC_43_out1_ready;
	wire phiC_43_out1_valid;

	wire sink_0_clk;
	wire sink_0_rst;
	wire [0 : 0]sink_0_in1_data;
	wire sink_0_in1_ready;
	wire sink_0_in1_valid;

	wire phi_7_clk;
	wire phi_7_rst;
	wire [0 : 0]phi_7_in1_data;
	wire phi_7_in1_ready;
	wire phi_7_in1_valid;
	wire [31 : 0]phi_7_in2_data;
	wire phi_7_in2_ready;
	wire phi_7_in2_valid;
	wire [31 : 0]phi_7_in3_data;
	wire phi_7_in3_ready;
	wire phi_7_in3_valid;
	wire [31 : 0]phi_7_out1_data;
	wire phi_7_out1_ready;
	wire phi_7_out1_valid;

	wire cst_3_clk;
	wire cst_3_rst;
	wire [0 : 0]cst_3_in1_data;
	wire cst_3_in1_ready;
	wire cst_3_in1_valid;
	wire [0 : 0]cst_3_out1_data;
	wire cst_3_out1_ready;
	wire cst_3_out1_valid;

	wire icmp_8_clk;
	wire icmp_8_rst;
	wire [31 : 0]icmp_8_in1_data;
	wire icmp_8_in1_ready;
	wire icmp_8_in1_valid;
	wire [31 : 0]icmp_8_in2_data;
	wire icmp_8_in2_ready;
	wire icmp_8_in2_valid;
	wire [0 : 0]icmp_8_out1_data;
	wire icmp_8_out1_ready;
	wire icmp_8_out1_valid;

	wire phi_n6_clk;
	wire phi_n6_rst;
	wire [31 : 0]phi_n6_in1_data;
	wire phi_n6_in1_ready;
	wire phi_n6_in1_valid;
	wire [31 : 0]phi_n6_in2_data;
	wire phi_n6_in2_ready;
	wire phi_n6_in2_valid;
	wire [31 : 0]phi_n6_out1_data;
	wire phi_n6_out1_ready;
	wire phi_n6_out1_valid;

	wire phi_n7_clk;
	wire phi_n7_rst;
	wire [2 : 0]phi_n7_in1_data;
	wire phi_n7_in1_ready;
	wire phi_n7_in1_valid;
	wire [2 : 0]phi_n7_in2_data;
	wire phi_n7_in2_ready;
	wire phi_n7_in2_valid;
	wire [2 : 0]phi_n7_out1_data;
	wire phi_n7_out1_ready;
	wire phi_n7_out1_valid;

	wire fork_1_clk;
	wire fork_1_rst;
	wire [31 : 0]fork_1_in1_data;
	wire fork_1_in1_ready;
	wire fork_1_in1_valid;
	wire [31 : 0]fork_1_out1_data;
	wire fork_1_out1_ready;
	wire fork_1_out1_valid;
	wire [31 : 0]fork_1_out2_data;
	wire fork_1_out2_ready;
	wire fork_1_out2_valid;

	wire branch_5_clk;
	wire branch_5_rst;
	wire [31 : 0]branch_5_in1_data;
	wire branch_5_in1_ready;
	wire branch_5_in1_valid;
	wire [0 : 0]branch_5_in2_data;
	wire branch_5_in2_ready;
	wire branch_5_in2_valid;
	wire [31 : 0]branch_5_out1_data;
	wire branch_5_out1_ready;
	wire branch_5_out1_valid;
	wire [31 : 0]branch_5_out2_data;
	wire branch_5_out2_ready;
	wire branch_5_out2_valid;

	wire branch_6_clk;
	wire branch_6_rst;
	wire [31 : 0]branch_6_in1_data;
	wire branch_6_in1_ready;
	wire branch_6_in1_valid;
	wire [0 : 0]branch_6_in2_data;
	wire branch_6_in2_ready;
	wire branch_6_in2_valid;
	wire [31 : 0]branch_6_out1_data;
	wire branch_6_out1_ready;
	wire branch_6_out1_valid;
	wire [31 : 0]branch_6_out2_data;
	wire branch_6_out2_ready;
	wire branch_6_out2_valid;

	wire branch_7_clk;
	wire branch_7_rst;
	wire [2 : 0]branch_7_in1_data;
	wire branch_7_in1_ready;
	wire branch_7_in1_valid;
	wire [0 : 0]branch_7_in2_data;
	wire branch_7_in2_ready;
	wire branch_7_in2_valid;
	wire [2 : 0]branch_7_out1_data;
	wire branch_7_out1_ready;
	wire branch_7_out1_valid;
	wire [2 : 0]branch_7_out2_data;
	wire branch_7_out2_ready;
	wire branch_7_out2_valid;

	wire fork_29_clk;
	wire fork_29_rst;
	wire [0 : 0]fork_29_in1_data;
	wire fork_29_in1_ready;
	wire fork_29_in1_valid;
	wire [0 : 0]fork_29_out1_data;
	wire fork_29_out1_ready;
	wire fork_29_out1_valid;
	wire [0 : 0]fork_29_out2_data;
	wire fork_29_out2_ready;
	wire fork_29_out2_valid;
	wire [0 : 0]fork_29_out3_data;
	wire fork_29_out3_ready;
	wire fork_29_out3_valid;
	wire [0 : 0]fork_29_out4_data;
	wire fork_29_out4_ready;
	wire fork_29_out4_valid;

	wire phiC_31_clk;
	wire phiC_31_rst;
	wire [0 : 0]phiC_31_in1_data;
	wire phiC_31_in1_ready;
	wire phiC_31_in1_valid;
	wire [0 : 0]phiC_31_in2_data;
	wire phiC_31_in2_ready;
	wire phiC_31_in2_valid;
	wire [0 : 0]phiC_31_out1_data;
	wire phiC_31_out1_ready;
	wire phiC_31_out1_valid;
	wire [0 : 0]phiC_31_out2_data;
	wire phiC_31_out2_ready;
	wire phiC_31_out2_valid;

	wire branchC_46_clk;
	wire branchC_46_rst;
	wire [0 : 0]branchC_46_in1_data;
	wire branchC_46_in1_ready;
	wire branchC_46_in1_valid;
	wire [0 : 0]branchC_46_in2_data;
	wire branchC_46_in2_ready;
	wire branchC_46_in2_valid;
	wire [0 : 0]branchC_46_out1_data;
	wire branchC_46_out1_ready;
	wire branchC_46_out1_valid;
	wire [0 : 0]branchC_46_out2_data;
	wire branchC_46_out2_ready;
	wire branchC_46_out2_valid;

	wire source_0_clk;
	wire source_0_rst;
	wire [0 : 0]source_0_out1_data;
	wire source_0_out1_ready;
	wire source_0_out1_valid;

	wire load_17_clk;
	wire load_17_rst;
	wire [31 : 0]load_17_in1_data;
	wire load_17_in1_ready;
	wire load_17_in1_valid;
	wire [2 : 0]load_17_in2_data;
	wire load_17_in2_ready;
	wire load_17_in2_valid;
	wire [31 : 0]load_17_out1_data;
	wire load_17_out1_ready;
	wire load_17_out1_valid;
	wire [2 : 0]load_17_out2_data;
	wire load_17_out2_ready;
	wire load_17_out2_valid;

	wire brCst_block5_clk;
	wire brCst_block5_rst;
	wire [0 : 0]brCst_block5_in1_data;
	wire brCst_block5_in1_ready;
	wire brCst_block5_in1_valid;
	wire [0 : 0]brCst_block5_out1_data;
	wire brCst_block5_out1_ready;
	wire brCst_block5_out1_valid;

	wire phi_n8_clk;
	wire phi_n8_rst;
	wire [2 : 0]phi_n8_in1_data;
	wire phi_n8_in1_ready;
	wire phi_n8_in1_valid;
	wire [2 : 0]phi_n8_out1_data;
	wire phi_n8_out1_ready;
	wire phi_n8_out1_valid;

	wire phi_n9_clk;
	wire phi_n9_rst;
	wire [31 : 0]phi_n9_in1_data;
	wire phi_n9_in1_ready;
	wire phi_n9_in1_valid;
	wire [31 : 0]phi_n9_out1_data;
	wire phi_n9_out1_ready;
	wire phi_n9_out1_valid;

	wire fork_16_clk;
	wire fork_16_rst;
	wire [2 : 0]fork_16_in1_data;
	wire fork_16_in1_ready;
	wire fork_16_in1_valid;
	wire [2 : 0]fork_16_out1_data;
	wire fork_16_out1_ready;
	wire fork_16_out1_valid;
	wire [2 : 0]fork_16_out2_data;
	wire fork_16_out2_ready;
	wire fork_16_out2_valid;

	wire branch_11_clk;
	wire branch_11_rst;
	wire [31 : 0]branch_11_in1_data;
	wire branch_11_in1_ready;
	wire branch_11_in1_valid;
	wire [0 : 0]branch_11_in2_data;
	wire branch_11_in2_ready;
	wire branch_11_in2_valid;
	wire [31 : 0]branch_11_out1_data;
	wire branch_11_out1_ready;
	wire branch_11_out1_valid;
	wire [31 : 0]branch_11_out2_data;
	wire branch_11_out2_ready;
	wire branch_11_out2_valid;

	wire branch_12_clk;
	wire branch_12_rst;
	wire [31 : 0]branch_12_in1_data;
	wire branch_12_in1_ready;
	wire branch_12_in1_valid;
	wire [0 : 0]branch_12_in2_data;
	wire branch_12_in2_ready;
	wire branch_12_in2_valid;
	wire [31 : 0]branch_12_out1_data;
	wire branch_12_out1_ready;
	wire branch_12_out1_valid;
	wire [31 : 0]branch_12_out2_data;
	wire branch_12_out2_ready;
	wire branch_12_out2_valid;

	wire branch_13_clk;
	wire branch_13_rst;
	wire [2 : 0]branch_13_in1_data;
	wire branch_13_in1_ready;
	wire branch_13_in1_valid;
	wire [0 : 0]branch_13_in2_data;
	wire branch_13_in2_ready;
	wire branch_13_in2_valid;
	wire [2 : 0]branch_13_out1_data;
	wire branch_13_out1_ready;
	wire branch_13_out1_valid;
	wire [2 : 0]branch_13_out2_data;
	wire branch_13_out2_ready;
	wire branch_13_out2_valid;

	wire fork_31_clk;
	wire fork_31_rst;
	wire [0 : 0]fork_31_in1_data;
	wire fork_31_in1_ready;
	wire fork_31_in1_valid;
	wire [0 : 0]fork_31_out1_data;
	wire fork_31_out1_ready;
	wire fork_31_out1_valid;
	wire [0 : 0]fork_31_out2_data;
	wire fork_31_out2_ready;
	wire fork_31_out2_valid;
	wire [0 : 0]fork_31_out3_data;
	wire fork_31_out3_ready;
	wire fork_31_out3_valid;
	wire [0 : 0]fork_31_out4_data;
	wire fork_31_out4_ready;
	wire fork_31_out4_valid;

	wire phiC_33_clk;
	wire phiC_33_rst;
	wire [0 : 0]phiC_33_in1_data;
	wire phiC_33_in1_ready;
	wire phiC_33_in1_valid;
	wire [0 : 0]phiC_33_out1_data;
	wire phiC_33_out1_ready;
	wire phiC_33_out1_valid;

	wire forkC_46_clk;
	wire forkC_46_rst;
	wire [0 : 0]forkC_46_in1_data;
	wire forkC_46_in1_ready;
	wire forkC_46_in1_valid;
	wire [0 : 0]forkC_46_out1_data;
	wire forkC_46_out1_ready;
	wire forkC_46_out1_valid;
	wire [0 : 0]forkC_46_out2_data;
	wire forkC_46_out2_ready;
	wire forkC_46_out2_valid;

	wire branchC_48_clk;
	wire branchC_48_rst;
	wire [0 : 0]branchC_48_in1_data;
	wire branchC_48_in1_ready;
	wire branchC_48_in1_valid;
	wire [0 : 0]branchC_48_in2_data;
	wire branchC_48_in2_ready;
	wire branchC_48_in2_valid;
	wire [0 : 0]branchC_48_out1_data;
	wire branchC_48_out1_ready;
	wire branchC_48_out1_valid;
	wire [0 : 0]branchC_48_out2_data;
	wire branchC_48_out2_ready;
	wire branchC_48_out2_valid;

	wire phi_38_clk;
	wire phi_38_rst;
	wire [0 : 0]phi_38_in1_data;
	wire phi_38_in1_ready;
	wire phi_38_in1_valid;
	wire [31 : 0]phi_38_in2_data;
	wire phi_38_in2_ready;
	wire phi_38_in2_valid;
	wire [31 : 0]phi_38_in3_data;
	wire phi_38_in3_ready;
	wire phi_38_in3_valid;
	wire [31 : 0]phi_38_out1_data;
	wire phi_38_out1_ready;
	wire phi_38_out1_valid;

	wire cst_9_clk;
	wire cst_9_rst;
	wire [0 : 0]cst_9_in1_data;
	wire cst_9_in1_ready;
	wire cst_9_in1_valid;
	wire [0 : 0]cst_9_out1_data;
	wire cst_9_out1_ready;
	wire cst_9_out1_valid;

	wire icmp_39_clk;
	wire icmp_39_rst;
	wire [31 : 0]icmp_39_in1_data;
	wire icmp_39_in1_ready;
	wire icmp_39_in1_valid;
	wire [31 : 0]icmp_39_in2_data;
	wire icmp_39_in2_ready;
	wire icmp_39_in2_valid;
	wire [0 : 0]icmp_39_out1_data;
	wire icmp_39_out1_ready;
	wire icmp_39_out1_valid;

	wire phi_n10_clk;
	wire phi_n10_rst;
	wire [31 : 0]phi_n10_in1_data;
	wire phi_n10_in1_ready;
	wire phi_n10_in1_valid;
	wire [31 : 0]phi_n10_in2_data;
	wire phi_n10_in2_ready;
	wire phi_n10_in2_valid;
	wire [31 : 0]phi_n10_out1_data;
	wire phi_n10_out1_ready;
	wire phi_n10_out1_valid;

	wire phi_n11_clk;
	wire phi_n11_rst;
	wire [31 : 0]phi_n11_in1_data;
	wire phi_n11_in1_ready;
	wire phi_n11_in1_valid;
	wire [31 : 0]phi_n11_in2_data;
	wire phi_n11_in2_ready;
	wire phi_n11_in2_valid;
	wire [31 : 0]phi_n11_out1_data;
	wire phi_n11_out1_ready;
	wire phi_n11_out1_valid;

	wire phi_n12_clk;
	wire phi_n12_rst;
	wire [9 : 0]phi_n12_in1_data;
	wire phi_n12_in1_ready;
	wire phi_n12_in1_valid;
	wire [9 : 0]phi_n12_in2_data;
	wire phi_n12_in2_ready;
	wire phi_n12_in2_valid;
	wire [9 : 0]phi_n12_out1_data;
	wire phi_n12_out1_ready;
	wire phi_n12_out1_valid;

	wire fork_5_clk;
	wire fork_5_rst;
	wire [31 : 0]fork_5_in1_data;
	wire fork_5_in1_ready;
	wire fork_5_in1_valid;
	wire [31 : 0]fork_5_out1_data;
	wire fork_5_out1_ready;
	wire fork_5_out1_valid;
	wire [31 : 0]fork_5_out2_data;
	wire fork_5_out2_ready;
	wire fork_5_out2_valid;

	wire branch_23_clk;
	wire branch_23_rst;
	wire [31 : 0]branch_23_in1_data;
	wire branch_23_in1_ready;
	wire branch_23_in1_valid;
	wire [0 : 0]branch_23_in2_data;
	wire branch_23_in2_ready;
	wire branch_23_in2_valid;
	wire [31 : 0]branch_23_out1_data;
	wire branch_23_out1_ready;
	wire branch_23_out1_valid;
	wire [31 : 0]branch_23_out2_data;
	wire branch_23_out2_ready;
	wire branch_23_out2_valid;

	wire branch_24_clk;
	wire branch_24_rst;
	wire [31 : 0]branch_24_in1_data;
	wire branch_24_in1_ready;
	wire branch_24_in1_valid;
	wire [0 : 0]branch_24_in2_data;
	wire branch_24_in2_ready;
	wire branch_24_in2_valid;
	wire [31 : 0]branch_24_out1_data;
	wire branch_24_out1_ready;
	wire branch_24_out1_valid;
	wire [31 : 0]branch_24_out2_data;
	wire branch_24_out2_ready;
	wire branch_24_out2_valid;

	wire branch_25_clk;
	wire branch_25_rst;
	wire [31 : 0]branch_25_in1_data;
	wire branch_25_in1_ready;
	wire branch_25_in1_valid;
	wire [0 : 0]branch_25_in2_data;
	wire branch_25_in2_ready;
	wire branch_25_in2_valid;
	wire [31 : 0]branch_25_out1_data;
	wire branch_25_out1_ready;
	wire branch_25_out1_valid;
	wire [31 : 0]branch_25_out2_data;
	wire branch_25_out2_ready;
	wire branch_25_out2_valid;

	wire branch_26_clk;
	wire branch_26_rst;
	wire [9 : 0]branch_26_in1_data;
	wire branch_26_in1_ready;
	wire branch_26_in1_valid;
	wire [0 : 0]branch_26_in2_data;
	wire branch_26_in2_ready;
	wire branch_26_in2_valid;
	wire [9 : 0]branch_26_out1_data;
	wire branch_26_out1_ready;
	wire branch_26_out1_valid;
	wire [9 : 0]branch_26_out2_data;
	wire branch_26_out2_ready;
	wire branch_26_out2_valid;

	wire fork_35_clk;
	wire fork_35_rst;
	wire [0 : 0]fork_35_in1_data;
	wire fork_35_in1_ready;
	wire fork_35_in1_valid;
	wire [0 : 0]fork_35_out1_data;
	wire fork_35_out1_ready;
	wire fork_35_out1_valid;
	wire [0 : 0]fork_35_out2_data;
	wire fork_35_out2_ready;
	wire fork_35_out2_valid;
	wire [0 : 0]fork_35_out3_data;
	wire fork_35_out3_ready;
	wire fork_35_out3_valid;
	wire [0 : 0]fork_35_out4_data;
	wire fork_35_out4_ready;
	wire fork_35_out4_valid;
	wire [0 : 0]fork_35_out5_data;
	wire fork_35_out5_ready;
	wire fork_35_out5_valid;

	wire phiC_37_clk;
	wire phiC_37_rst;
	wire [0 : 0]phiC_37_in1_data;
	wire phiC_37_in1_ready;
	wire phiC_37_in1_valid;
	wire [0 : 0]phiC_37_in2_data;
	wire phiC_37_in2_ready;
	wire phiC_37_in2_valid;
	wire [0 : 0]phiC_37_out1_data;
	wire phiC_37_out1_ready;
	wire phiC_37_out1_valid;
	wire [0 : 0]phiC_37_out2_data;
	wire phiC_37_out2_ready;
	wire phiC_37_out2_valid;

	wire branchC_52_clk;
	wire branchC_52_rst;
	wire [0 : 0]branchC_52_in1_data;
	wire branchC_52_in1_ready;
	wire branchC_52_in1_valid;
	wire [0 : 0]branchC_52_in2_data;
	wire branchC_52_in2_ready;
	wire branchC_52_in2_valid;
	wire [0 : 0]branchC_52_out1_data;
	wire branchC_52_out1_ready;
	wire branchC_52_out1_valid;
	wire [0 : 0]branchC_52_out2_data;
	wire branchC_52_out2_ready;
	wire branchC_52_out2_valid;

	wire source_3_clk;
	wire source_3_rst;
	wire [0 : 0]source_3_out1_data;
	wire source_3_out1_ready;
	wire source_3_out1_valid;

	wire load_21_clk;
	wire load_21_rst;
	wire [31 : 0]load_21_in1_data;
	wire load_21_in1_ready;
	wire load_21_in1_valid;
	wire [31 : 0]load_21_in2_data;
	wire load_21_in2_ready;
	wire load_21_in2_valid;
	wire [31 : 0]load_21_out1_data;
	wire load_21_out1_ready;
	wire load_21_out1_valid;
	wire [31 : 0]load_21_out2_data;
	wire load_21_out2_ready;
	wire load_21_out2_valid;

	wire icmp_22_clk;
	wire icmp_22_rst;
	wire [31 : 0]icmp_22_in1_data;
	wire icmp_22_in1_ready;
	wire icmp_22_in1_valid;
	wire [31 : 0]icmp_22_in2_data;
	wire icmp_22_in2_ready;
	wire icmp_22_in2_valid;
	wire [0 : 0]icmp_22_out1_data;
	wire icmp_22_out1_ready;
	wire icmp_22_out1_valid;

	wire zext_23_clk;
	wire zext_23_rst;
	wire [0 : 0]zext_23_in1_data;
	wire zext_23_in1_ready;
	wire zext_23_in1_valid;
	wire [0 : 0]zext_23_out1_data;
	wire zext_23_out1_ready;
	wire zext_23_out1_valid;

	wire add_24_clk;
	wire add_24_rst;
	wire [31 : 0]add_24_in1_data;
	wire add_24_in1_ready;
	wire add_24_in1_valid;
	wire [31 : 0]add_24_in2_data;
	wire add_24_in2_ready;
	wire add_24_in2_valid;
	wire [31 : 0]add_24_out1_data;
	wire add_24_out1_ready;
	wire add_24_out1_valid;

	wire store_1_clk;
	wire store_1_rst;
	wire [31 : 0]store_1_in1_data;
	wire store_1_in1_ready;
	wire store_1_in1_valid;
	wire [2 : 0]store_1_in2_data;
	wire store_1_in2_ready;
	wire store_1_in2_valid;
	wire [31 : 0]store_1_out1_data;
	wire store_1_out1_ready;
	wire store_1_out1_valid;
	wire [2 : 0]store_1_out2_data;
	wire store_1_out2_ready;
	wire store_1_out2_valid;

	wire cst_4_clk;
	wire cst_4_rst;
	wire [0 : 0]cst_4_in1_data;
	wire cst_4_in1_ready;
	wire cst_4_in1_valid;
	wire [0 : 0]cst_4_out1_data;
	wire cst_4_out1_ready;
	wire cst_4_out1_valid;

	wire add_27_clk;
	wire add_27_rst;
	wire [2 : 0]add_27_in1_data;
	wire add_27_in1_ready;
	wire add_27_in1_valid;
	wire [2 : 0]add_27_in2_data;
	wire add_27_in2_ready;
	wire add_27_in2_valid;
	wire [2 : 0]add_27_out1_data;
	wire add_27_out1_ready;
	wire add_27_out1_valid;

	wire cst_5_clk;
	wire cst_5_rst;
	wire [2 : 0]cst_5_in1_data;
	wire cst_5_in1_ready;
	wire cst_5_in1_valid;
	wire [2 : 0]cst_5_out1_data;
	wire cst_5_out1_ready;
	wire cst_5_out1_valid;

	wire icmp_28_clk;
	wire icmp_28_rst;
	wire [2 : 0]icmp_28_in1_data;
	wire icmp_28_in1_ready;
	wire icmp_28_in1_valid;
	wire [2 : 0]icmp_28_in2_data;
	wire icmp_28_in2_ready;
	wire icmp_28_in2_valid;
	wire [0 : 0]icmp_28_out1_data;
	wire icmp_28_out1_ready;
	wire icmp_28_out1_valid;

	wire phi_n3_clk;
	wire phi_n3_rst;
	wire [31 : 0]phi_n3_in1_data;
	wire phi_n3_in1_ready;
	wire phi_n3_in1_valid;
	wire [31 : 0]phi_n3_in2_data;
	wire phi_n3_in2_ready;
	wire phi_n3_in2_valid;
	wire [31 : 0]phi_n3_out1_data;
	wire phi_n3_out1_ready;
	wire phi_n3_out1_valid;

	wire phi_n4_clk;
	wire phi_n4_rst;
	wire [31 : 0]phi_n4_in1_data;
	wire phi_n4_in1_ready;
	wire phi_n4_in1_valid;
	wire [31 : 0]phi_n4_in2_data;
	wire phi_n4_in2_ready;
	wire phi_n4_in2_valid;
	wire [31 : 0]phi_n4_out1_data;
	wire phi_n4_out1_ready;
	wire phi_n4_out1_valid;

	wire phi_n5_clk;
	wire phi_n5_rst;
	wire [2 : 0]phi_n5_in1_data;
	wire phi_n5_in1_ready;
	wire phi_n5_in1_valid;
	wire [2 : 0]phi_n5_in2_data;
	wire phi_n5_in2_ready;
	wire phi_n5_in2_valid;
	wire [2 : 0]phi_n5_out1_data;
	wire phi_n5_out1_ready;
	wire phi_n5_out1_valid;

	wire fork_2_clk;
	wire fork_2_rst;
	wire [31 : 0]fork_2_in1_data;
	wire fork_2_in1_ready;
	wire fork_2_in1_valid;
	wire [31 : 0]fork_2_out1_data;
	wire fork_2_out1_ready;
	wire fork_2_out1_valid;
	wire [31 : 0]fork_2_out2_data;
	wire fork_2_out2_ready;
	wire fork_2_out2_valid;

	wire fork_3_clk;
	wire fork_3_rst;
	wire [2 : 0]fork_3_in1_data;
	wire fork_3_in1_ready;
	wire fork_3_in1_valid;
	wire [2 : 0]fork_3_out1_data;
	wire fork_3_out1_ready;
	wire fork_3_out1_valid;
	wire [2 : 0]fork_3_out2_data;
	wire fork_3_out2_ready;
	wire fork_3_out2_valid;

	wire fork_12_clk;
	wire fork_12_rst;
	wire [31 : 0]fork_12_in1_data;
	wire fork_12_in1_ready;
	wire fork_12_in1_valid;
	wire [31 : 0]fork_12_out1_data;
	wire fork_12_out1_ready;
	wire fork_12_out1_valid;
	wire [31 : 0]fork_12_out2_data;
	wire fork_12_out2_ready;
	wire fork_12_out2_valid;

	wire fork_13_clk;
	wire fork_13_rst;
	wire [2 : 0]fork_13_in1_data;
	wire fork_13_in1_ready;
	wire fork_13_in1_valid;
	wire [2 : 0]fork_13_out1_data;
	wire fork_13_out1_ready;
	wire fork_13_out1_valid;
	wire [2 : 0]fork_13_out2_data;
	wire fork_13_out2_ready;
	wire fork_13_out2_valid;

	wire branch_14_clk;
	wire branch_14_rst;
	wire [31 : 0]branch_14_in1_data;
	wire branch_14_in1_ready;
	wire branch_14_in1_valid;
	wire [0 : 0]branch_14_in2_data;
	wire branch_14_in2_ready;
	wire branch_14_in2_valid;
	wire [31 : 0]branch_14_out1_data;
	wire branch_14_out1_ready;
	wire branch_14_out1_valid;
	wire [31 : 0]branch_14_out2_data;
	wire branch_14_out2_ready;
	wire branch_14_out2_valid;

	wire branch_15_clk;
	wire branch_15_rst;
	wire [2 : 0]branch_15_in1_data;
	wire branch_15_in1_ready;
	wire branch_15_in1_valid;
	wire [0 : 0]branch_15_in2_data;
	wire branch_15_in2_ready;
	wire branch_15_in2_valid;
	wire [2 : 0]branch_15_out1_data;
	wire branch_15_out1_ready;
	wire branch_15_out1_valid;
	wire [2 : 0]branch_15_out2_data;
	wire branch_15_out2_ready;
	wire branch_15_out2_valid;

	wire fork_32_clk;
	wire fork_32_rst;
	wire [0 : 0]fork_32_in1_data;
	wire fork_32_in1_ready;
	wire fork_32_in1_valid;
	wire [0 : 0]fork_32_out1_data;
	wire fork_32_out1_ready;
	wire fork_32_out1_valid;
	wire [0 : 0]fork_32_out2_data;
	wire fork_32_out2_ready;
	wire fork_32_out2_valid;
	wire [0 : 0]fork_32_out3_data;
	wire fork_32_out3_ready;
	wire fork_32_out3_valid;

	wire cst_17_clk;
	wire cst_17_rst;
	wire [0 : 0]cst_17_in1_data;
	wire cst_17_in1_ready;
	wire cst_17_in1_valid;
	wire [0 : 0]cst_17_out1_data;
	wire cst_17_out1_ready;
	wire cst_17_out1_valid;

	wire phiC_34_clk;
	wire phiC_34_rst;
	wire [0 : 0]phiC_34_in1_data;
	wire phiC_34_in1_ready;
	wire phiC_34_in1_valid;
	wire [0 : 0]phiC_34_in2_data;
	wire phiC_34_in2_ready;
	wire phiC_34_in2_valid;
	wire [0 : 0]phiC_34_out1_data;
	wire phiC_34_out1_ready;
	wire phiC_34_out1_valid;

	wire forkC_47_clk;
	wire forkC_47_rst;
	wire [0 : 0]forkC_47_in1_data;
	wire forkC_47_in1_ready;
	wire forkC_47_in1_valid;
	wire [0 : 0]forkC_47_out1_data;
	wire forkC_47_out1_ready;
	wire forkC_47_out1_valid;
	wire [0 : 0]forkC_47_out2_data;
	wire forkC_47_out2_ready;
	wire forkC_47_out2_valid;

	wire branchC_49_clk;
	wire branchC_49_rst;
	wire [0 : 0]branchC_49_in1_data;
	wire branchC_49_in1_ready;
	wire branchC_49_in1_valid;
	wire [0 : 0]branchC_49_in2_data;
	wire branchC_49_in2_ready;
	wire branchC_49_in2_valid;
	wire [0 : 0]branchC_49_out1_data;
	wire branchC_49_out1_ready;
	wire branchC_49_out1_valid;
	wire [0 : 0]branchC_49_out2_data;
	wire branchC_49_out2_ready;
	wire branchC_49_out2_valid;

	wire source_1_clk;
	wire source_1_rst;
	wire [0 : 0]source_1_out1_data;
	wire source_1_out1_ready;
	wire source_1_out1_valid;

	wire source_2_clk;
	wire source_2_rst;
	wire [2 : 0]source_2_out1_data;
	wire source_2_out1_ready;
	wire source_2_out1_valid;

	wire load_12_clk;
	wire load_12_rst;
	wire [31 : 0]load_12_in1_data;
	wire load_12_in1_ready;
	wire load_12_in1_valid;
	wire [31 : 0]load_12_in2_data;
	wire load_12_in2_ready;
	wire load_12_in2_valid;
	wire [31 : 0]load_12_out1_data;
	wire load_12_out1_ready;
	wire load_12_out1_valid;
	wire [31 : 0]load_12_out2_data;
	wire load_12_out2_ready;
	wire load_12_out2_valid;

	wire icmp_13_clk;
	wire icmp_13_rst;
	wire [31 : 0]icmp_13_in1_data;
	wire icmp_13_in1_ready;
	wire icmp_13_in1_valid;
	wire [31 : 0]icmp_13_in2_data;
	wire icmp_13_in2_ready;
	wire icmp_13_in2_valid;
	wire [0 : 0]icmp_13_out1_data;
	wire icmp_13_out1_ready;
	wire icmp_13_out1_valid;

	wire phi_n0_clk;
	wire phi_n0_rst;
	wire [31 : 0]phi_n0_in1_data;
	wire phi_n0_in1_ready;
	wire phi_n0_in1_valid;
	wire [31 : 0]phi_n0_out1_data;
	wire phi_n0_out1_ready;
	wire phi_n0_out1_valid;

	wire phi_n1_clk;
	wire phi_n1_rst;
	wire [31 : 0]phi_n1_in1_data;
	wire phi_n1_in1_ready;
	wire phi_n1_in1_valid;
	wire [31 : 0]phi_n1_out1_data;
	wire phi_n1_out1_ready;
	wire phi_n1_out1_valid;

	wire phi_n2_clk;
	wire phi_n2_rst;
	wire [2 : 0]phi_n2_in1_data;
	wire phi_n2_in1_ready;
	wire phi_n2_in1_valid;
	wire [2 : 0]phi_n2_out1_data;
	wire phi_n2_out1_ready;
	wire phi_n2_out1_valid;

	wire fork_9_clk;
	wire fork_9_rst;
	wire [31 : 0]fork_9_in1_data;
	wire fork_9_in1_ready;
	wire fork_9_in1_valid;
	wire [31 : 0]fork_9_out1_data;
	wire fork_9_out1_ready;
	wire fork_9_out1_valid;
	wire [31 : 0]fork_9_out2_data;
	wire fork_9_out2_ready;
	wire fork_9_out2_valid;

	wire fork_10_clk;
	wire fork_10_rst;
	wire [31 : 0]fork_10_in1_data;
	wire fork_10_in1_ready;
	wire fork_10_in1_valid;
	wire [31 : 0]fork_10_out1_data;
	wire fork_10_out1_ready;
	wire fork_10_out1_valid;
	wire [31 : 0]fork_10_out2_data;
	wire fork_10_out2_ready;
	wire fork_10_out2_valid;

	wire branch_8_clk;
	wire branch_8_rst;
	wire [31 : 0]branch_8_in1_data;
	wire branch_8_in1_ready;
	wire branch_8_in1_valid;
	wire [0 : 0]branch_8_in2_data;
	wire branch_8_in2_ready;
	wire branch_8_in2_valid;
	wire [31 : 0]branch_8_out1_data;
	wire branch_8_out1_ready;
	wire branch_8_out1_valid;
	wire [31 : 0]branch_8_out2_data;
	wire branch_8_out2_ready;
	wire branch_8_out2_valid;

	wire branch_9_clk;
	wire branch_9_rst;
	wire [31 : 0]branch_9_in1_data;
	wire branch_9_in1_ready;
	wire branch_9_in1_valid;
	wire [0 : 0]branch_9_in2_data;
	wire branch_9_in2_ready;
	wire branch_9_in2_valid;
	wire [31 : 0]branch_9_out1_data;
	wire branch_9_out1_ready;
	wire branch_9_out1_valid;
	wire [31 : 0]branch_9_out2_data;
	wire branch_9_out2_ready;
	wire branch_9_out2_valid;

	wire branch_10_clk;
	wire branch_10_rst;
	wire [2 : 0]branch_10_in1_data;
	wire branch_10_in1_ready;
	wire branch_10_in1_valid;
	wire [0 : 0]branch_10_in2_data;
	wire branch_10_in2_ready;
	wire branch_10_in2_valid;
	wire [2 : 0]branch_10_out1_data;
	wire branch_10_out1_ready;
	wire branch_10_out1_valid;
	wire [2 : 0]branch_10_out2_data;
	wire branch_10_out2_ready;
	wire branch_10_out2_valid;

	wire fork_30_clk;
	wire fork_30_rst;
	wire [0 : 0]fork_30_in1_data;
	wire fork_30_in1_ready;
	wire fork_30_in1_valid;
	wire [0 : 0]fork_30_out1_data;
	wire fork_30_out1_ready;
	wire fork_30_out1_valid;
	wire [0 : 0]fork_30_out2_data;
	wire fork_30_out2_ready;
	wire fork_30_out2_valid;
	wire [0 : 0]fork_30_out3_data;
	wire fork_30_out3_ready;
	wire fork_30_out3_valid;
	wire [0 : 0]fork_30_out4_data;
	wire fork_30_out4_ready;
	wire fork_30_out4_valid;

	wire phiC_32_clk;
	wire phiC_32_rst;
	wire [0 : 0]phiC_32_in1_data;
	wire phiC_32_in1_ready;
	wire phiC_32_in1_valid;
	wire [0 : 0]phiC_32_out1_data;
	wire phiC_32_out1_ready;
	wire phiC_32_out1_valid;

	wire branchC_47_clk;
	wire branchC_47_rst;
	wire [0 : 0]branchC_47_in1_data;
	wire branchC_47_in1_ready;
	wire branchC_47_in1_valid;
	wire [0 : 0]branchC_47_in2_data;
	wire branchC_47_in2_ready;
	wire branchC_47_in2_valid;
	wire [0 : 0]branchC_47_out1_data;
	wire branchC_47_out1_ready;
	wire branchC_47_out1_valid;
	wire [0 : 0]branchC_47_out2_data;
	wire branchC_47_out2_ready;
	wire branchC_47_out2_valid;

	wire phi_64_clk;
	wire phi_64_rst;
	wire [0 : 0]phi_64_in1_data;
	wire phi_64_in1_ready;
	wire phi_64_in1_valid;
	wire [31 : 0]phi_64_in2_data;
	wire phi_64_in2_ready;
	wire phi_64_in2_valid;
	wire [31 : 0]phi_64_in3_data;
	wire phi_64_in3_ready;
	wire phi_64_in3_valid;
	wire [31 : 0]phi_64_out1_data;
	wire phi_64_out1_ready;
	wire phi_64_out1_valid;

	wire phi_65_clk;
	wire phi_65_rst;
	wire [0 : 0]phi_65_in1_data;
	wire phi_65_in1_ready;
	wire phi_65_in1_valid;
	wire [31 : 0]phi_65_in2_data;
	wire phi_65_in2_ready;
	wire phi_65_in2_valid;
	wire [31 : 0]phi_65_in3_data;
	wire phi_65_in3_ready;
	wire phi_65_in3_valid;
	wire [31 : 0]phi_65_out1_data;
	wire phi_65_out1_ready;
	wire phi_65_out1_valid;

	wire cst_13_clk;
	wire cst_13_rst;
	wire [0 : 0]cst_13_in1_data;
	wire cst_13_in1_ready;
	wire cst_13_in1_valid;
	wire [0 : 0]cst_13_out1_data;
	wire cst_13_out1_ready;
	wire cst_13_out1_valid;

	wire add_66_clk;
	wire add_66_rst;
	wire [9 : 0]add_66_in1_data;
	wire add_66_in1_ready;
	wire add_66_in1_valid;
	wire [9 : 0]add_66_in2_data;
	wire add_66_in2_ready;
	wire add_66_in2_valid;
	wire [9 : 0]add_66_out1_data;
	wire add_66_out1_ready;
	wire add_66_out1_valid;

	wire cst_14_clk;
	wire cst_14_rst;
	wire [9 : 0]cst_14_in1_data;
	wire cst_14_in1_ready;
	wire cst_14_in1_valid;
	wire [9 : 0]cst_14_out1_data;
	wire cst_14_out1_ready;
	wire cst_14_out1_valid;

	wire icmp_67_clk;
	wire icmp_67_rst;
	wire [9 : 0]icmp_67_in1_data;
	wire icmp_67_in1_ready;
	wire icmp_67_in1_valid;
	wire [9 : 0]icmp_67_in2_data;
	wire icmp_67_in2_ready;
	wire icmp_67_in2_valid;
	wire [0 : 0]icmp_67_out1_data;
	wire icmp_67_out1_ready;
	wire icmp_67_out1_valid;

	wire phi_n16_clk;
	wire phi_n16_rst;
	wire [9 : 0]phi_n16_in1_data;
	wire phi_n16_in1_ready;
	wire phi_n16_in1_valid;
	wire [9 : 0]phi_n16_in2_data;
	wire phi_n16_in2_ready;
	wire phi_n16_in2_valid;
	wire [9 : 0]phi_n16_out1_data;
	wire phi_n16_out1_ready;
	wire phi_n16_out1_valid;

	wire fork_8_clk;
	wire fork_8_rst;
	wire [9 : 0]fork_8_in1_data;
	wire fork_8_in1_ready;
	wire fork_8_in1_valid;
	wire [9 : 0]fork_8_out1_data;
	wire fork_8_out1_ready;
	wire fork_8_out1_valid;
	wire [9 : 0]fork_8_out2_data;
	wire fork_8_out2_ready;
	wire fork_8_out2_valid;

	wire branch_41_clk;
	wire branch_41_rst;
	wire [31 : 0]branch_41_in1_data;
	wire branch_41_in1_ready;
	wire branch_41_in1_valid;
	wire [0 : 0]branch_41_in2_data;
	wire branch_41_in2_ready;
	wire branch_41_in2_valid;
	wire [31 : 0]branch_41_out1_data;
	wire branch_41_out1_ready;
	wire branch_41_out1_valid;
	wire [31 : 0]branch_41_out2_data;
	wire branch_41_out2_ready;
	wire branch_41_out2_valid;

	wire branch_42_clk;
	wire branch_42_rst;
	wire [31 : 0]branch_42_in1_data;
	wire branch_42_in1_ready;
	wire branch_42_in1_valid;
	wire [0 : 0]branch_42_in2_data;
	wire branch_42_in2_ready;
	wire branch_42_in2_valid;
	wire [31 : 0]branch_42_out1_data;
	wire branch_42_out1_ready;
	wire branch_42_out1_valid;
	wire [31 : 0]branch_42_out2_data;
	wire branch_42_out2_ready;
	wire branch_42_out2_valid;

	wire branch_43_clk;
	wire branch_43_rst;
	wire [9 : 0]branch_43_in1_data;
	wire branch_43_in1_ready;
	wire branch_43_in1_valid;
	wire [0 : 0]branch_43_in2_data;
	wire branch_43_in2_ready;
	wire branch_43_in2_valid;
	wire [9 : 0]branch_43_out1_data;
	wire branch_43_out1_ready;
	wire branch_43_out1_valid;
	wire [9 : 0]branch_43_out2_data;
	wire branch_43_out2_ready;
	wire branch_43_out2_valid;

	wire fork_40_clk;
	wire fork_40_rst;
	wire [0 : 0]fork_40_in1_data;
	wire fork_40_in1_ready;
	wire fork_40_in1_valid;
	wire [0 : 0]fork_40_out1_data;
	wire fork_40_out1_ready;
	wire fork_40_out1_valid;
	wire [0 : 0]fork_40_out2_data;
	wire fork_40_out2_ready;
	wire fork_40_out2_valid;
	wire [0 : 0]fork_40_out3_data;
	wire fork_40_out3_ready;
	wire fork_40_out3_valid;
	wire [0 : 0]fork_40_out4_data;
	wire fork_40_out4_ready;
	wire fork_40_out4_valid;

	wire phiC_42_clk;
	wire phiC_42_rst;
	wire [0 : 0]phiC_42_in1_data;
	wire phiC_42_in1_ready;
	wire phiC_42_in1_valid;
	wire [0 : 0]phiC_42_in2_data;
	wire phiC_42_in2_ready;
	wire phiC_42_in2_valid;
	wire [0 : 0]phiC_42_out1_data;
	wire phiC_42_out1_ready;
	wire phiC_42_out1_valid;
	wire [0 : 0]phiC_42_out2_data;
	wire phiC_42_out2_ready;
	wire phiC_42_out2_valid;

	wire branchC_57_clk;
	wire branchC_57_rst;
	wire [0 : 0]branchC_57_in1_data;
	wire branchC_57_in1_ready;
	wire branchC_57_in1_valid;
	wire [0 : 0]branchC_57_in2_data;
	wire branchC_57_in2_ready;
	wire branchC_57_in2_valid;
	wire [0 : 0]branchC_57_out1_data;
	wire branchC_57_out1_ready;
	wire branchC_57_out1_valid;
	wire [0 : 0]branchC_57_out2_data;
	wire branchC_57_out2_ready;
	wire branchC_57_out2_valid;

	wire source_7_clk;
	wire source_7_rst;
	wire [0 : 0]source_7_out1_data;
	wire source_7_out1_ready;
	wire source_7_out1_valid;

	wire source_8_clk;
	wire source_8_rst;
	wire [9 : 0]source_8_out1_data;
	wire source_8_out1_ready;
	wire source_8_out1_valid;

	wire fork_61_clk;
	wire fork_61_rst;
	wire [0 : 0]fork_61_in1_data;
	wire fork_61_in1_ready;
	wire fork_61_in1_valid;
	wire [0 : 0]fork_61_out1_data;
	wire fork_61_out1_ready;
	wire fork_61_out1_valid;
	wire [0 : 0]fork_61_out2_data;
	wire fork_61_out2_ready;
	wire fork_61_out2_valid;

	wire cst_11_clk;
	wire cst_11_rst;
	wire [0 : 0]cst_11_in1_data;
	wire cst_11_in1_ready;
	wire cst_11_in1_valid;
	wire [0 : 0]cst_11_out1_data;
	wire cst_11_out1_ready;
	wire cst_11_out1_valid;

	wire add_58_clk;
	wire add_58_rst;
	wire [31 : 0]add_58_in1_data;
	wire add_58_in1_ready;
	wire add_58_in1_valid;
	wire [31 : 0]add_58_in2_data;
	wire add_58_in2_ready;
	wire add_58_in2_valid;
	wire [31 : 0]add_58_out1_data;
	wire add_58_out1_ready;
	wire add_58_out1_valid;

	wire cst_12_clk;
	wire cst_12_rst;
	wire [31 : 0]cst_12_in1_data;
	wire cst_12_in1_ready;
	wire cst_12_in1_valid;
	wire [31 : 0]cst_12_out1_data;
	wire cst_12_out1_ready;
	wire cst_12_out1_valid;

	wire add_59_clk;
	wire add_59_rst;
	wire [31 : 0]add_59_in1_data;
	wire add_59_in1_ready;
	wire add_59_in1_valid;
	wire [31 : 0]add_59_in2_data;
	wire add_59_in2_ready;
	wire add_59_in2_valid;
	wire [31 : 0]add_59_out1_data;
	wire add_59_out1_ready;
	wire add_59_out1_valid;

	wire load_62_clk;
	wire load_62_rst;
	wire [31 : 0]load_62_in1_data;
	wire load_62_in1_ready;
	wire load_62_in1_valid;
	wire [31 : 0]load_62_in2_data;
	wire load_62_in2_ready;
	wire load_62_in2_valid;
	wire [31 : 0]load_62_out1_data;
	wire load_62_out1_ready;
	wire load_62_out1_valid;
	wire [31 : 0]load_62_out2_data;
	wire load_62_out2_ready;
	wire load_62_out2_valid;

	wire brCst_block13_clk;
	wire brCst_block13_rst;
	wire [0 : 0]brCst_block13_in1_data;
	wire brCst_block13_in1_ready;
	wire brCst_block13_in1_valid;
	wire [0 : 0]brCst_block13_out1_data;
	wire brCst_block13_out1_ready;
	wire brCst_block13_out1_valid;

	wire phi_n13_clk;
	wire phi_n13_rst;
	wire [31 : 0]phi_n13_in1_data;
	wire phi_n13_in1_ready;
	wire phi_n13_in1_valid;
	wire [31 : 0]phi_n13_out1_data;
	wire phi_n13_out1_ready;
	wire phi_n13_out1_valid;

	wire phi_n14_clk;
	wire phi_n14_rst;
	wire [31 : 0]phi_n14_in1_data;
	wire phi_n14_in1_ready;
	wire phi_n14_in1_valid;
	wire [31 : 0]phi_n14_out1_data;
	wire phi_n14_out1_ready;
	wire phi_n14_out1_valid;

	wire phi_n15_clk;
	wire phi_n15_rst;
	wire [9 : 0]phi_n15_in1_data;
	wire phi_n15_in1_ready;
	wire phi_n15_in1_valid;
	wire [9 : 0]phi_n15_out1_data;
	wire phi_n15_out1_ready;
	wire phi_n15_out1_valid;

	wire branch_38_clk;
	wire branch_38_rst;
	wire [31 : 0]branch_38_in1_data;
	wire branch_38_in1_ready;
	wire branch_38_in1_valid;
	wire [0 : 0]branch_38_in2_data;
	wire branch_38_in2_ready;
	wire branch_38_in2_valid;
	wire [31 : 0]branch_38_out1_data;
	wire branch_38_out1_ready;
	wire branch_38_out1_valid;
	wire [31 : 0]branch_38_out2_data;
	wire branch_38_out2_ready;
	wire branch_38_out2_valid;

	wire branch_39_clk;
	wire branch_39_rst;
	wire [31 : 0]branch_39_in1_data;
	wire branch_39_in1_ready;
	wire branch_39_in1_valid;
	wire [0 : 0]branch_39_in2_data;
	wire branch_39_in2_ready;
	wire branch_39_in2_valid;
	wire [31 : 0]branch_39_out1_data;
	wire branch_39_out1_ready;
	wire branch_39_out1_valid;
	wire [31 : 0]branch_39_out2_data;
	wire branch_39_out2_ready;
	wire branch_39_out2_valid;

	wire branch_40_clk;
	wire branch_40_rst;
	wire [9 : 0]branch_40_in1_data;
	wire branch_40_in1_ready;
	wire branch_40_in1_valid;
	wire [0 : 0]branch_40_in2_data;
	wire branch_40_in2_ready;
	wire branch_40_in2_valid;
	wire [9 : 0]branch_40_out1_data;
	wire branch_40_out1_ready;
	wire branch_40_out1_valid;
	wire [9 : 0]branch_40_out2_data;
	wire branch_40_out2_ready;
	wire branch_40_out2_valid;

	wire fork_39_clk;
	wire fork_39_rst;
	wire [0 : 0]fork_39_in1_data;
	wire fork_39_in1_ready;
	wire fork_39_in1_valid;
	wire [0 : 0]fork_39_out1_data;
	wire fork_39_out1_ready;
	wire fork_39_out1_valid;
	wire [0 : 0]fork_39_out2_data;
	wire fork_39_out2_ready;
	wire fork_39_out2_valid;
	wire [0 : 0]fork_39_out3_data;
	wire fork_39_out3_ready;
	wire fork_39_out3_valid;
	wire [0 : 0]fork_39_out4_data;
	wire fork_39_out4_ready;
	wire fork_39_out4_valid;

	wire phiC_41_clk;
	wire phiC_41_rst;
	wire [0 : 0]phiC_41_in1_data;
	wire phiC_41_in1_ready;
	wire phiC_41_in1_valid;
	wire [0 : 0]phiC_41_out1_data;
	wire phiC_41_out1_ready;
	wire phiC_41_out1_valid;

	wire forkC_54_clk;
	wire forkC_54_rst;
	wire [0 : 0]forkC_54_in1_data;
	wire forkC_54_in1_ready;
	wire forkC_54_in1_valid;
	wire [0 : 0]forkC_54_out1_data;
	wire forkC_54_out1_ready;
	wire forkC_54_out1_valid;
	wire [0 : 0]forkC_54_out2_data;
	wire forkC_54_out2_ready;
	wire forkC_54_out2_valid;

	wire branchC_56_clk;
	wire branchC_56_rst;
	wire [0 : 0]branchC_56_in1_data;
	wire branchC_56_in1_ready;
	wire branchC_56_in1_valid;
	wire [0 : 0]branchC_56_in2_data;
	wire branchC_56_in2_ready;
	wire branchC_56_in2_valid;
	wire [0 : 0]branchC_56_out1_data;
	wire branchC_56_out1_ready;
	wire branchC_56_out1_valid;
	wire [0 : 0]branchC_56_out2_data;
	wire branchC_56_out2_ready;
	wire branchC_56_out2_valid;

	wire source_5_clk;
	wire source_5_rst;
	wire [0 : 0]source_5_out1_data;
	wire source_5_out1_ready;
	wire source_5_out1_valid;

	wire source_6_clk;
	wire source_6_rst;
	wire [31 : 0]source_6_out1_data;
	wire source_6_out1_ready;
	wire source_6_out1_valid;

	wire load_43_clk;
	wire load_43_rst;
	wire [31 : 0]load_43_in1_data;
	wire load_43_in1_ready;
	wire load_43_in1_valid;
	wire [31 : 0]load_43_in2_data;
	wire load_43_in2_ready;
	wire load_43_in2_valid;
	wire [31 : 0]load_43_out1_data;
	wire load_43_out1_ready;
	wire load_43_out1_valid;
	wire [31 : 0]load_43_out2_data;
	wire load_43_out2_ready;
	wire load_43_out2_valid;

	wire icmp_44_clk;
	wire icmp_44_rst;
	wire [31 : 0]icmp_44_in1_data;
	wire icmp_44_in1_ready;
	wire icmp_44_in1_valid;
	wire [31 : 0]icmp_44_in2_data;
	wire icmp_44_in2_ready;
	wire icmp_44_in2_valid;
	wire [0 : 0]icmp_44_out1_data;
	wire icmp_44_out1_ready;
	wire icmp_44_out1_valid;

	wire phi_n21_clk;
	wire phi_n21_rst;
	wire [31 : 0]phi_n21_in1_data;
	wire phi_n21_in1_ready;
	wire phi_n21_in1_valid;
	wire [31 : 0]phi_n21_out1_data;
	wire phi_n21_out1_ready;
	wire phi_n21_out1_valid;

	wire phi_n22_clk;
	wire phi_n22_rst;
	wire [31 : 0]phi_n22_in1_data;
	wire phi_n22_in1_ready;
	wire phi_n22_in1_valid;
	wire [31 : 0]phi_n22_out1_data;
	wire phi_n22_out1_ready;
	wire phi_n22_out1_valid;

	wire phi_n23_clk;
	wire phi_n23_rst;
	wire [31 : 0]phi_n23_in1_data;
	wire phi_n23_in1_ready;
	wire phi_n23_in1_valid;
	wire [31 : 0]phi_n23_out1_data;
	wire phi_n23_out1_ready;
	wire phi_n23_out1_valid;

	wire phi_n24_clk;
	wire phi_n24_rst;
	wire [9 : 0]phi_n24_in1_data;
	wire phi_n24_in1_ready;
	wire phi_n24_in1_valid;
	wire [9 : 0]phi_n24_out1_data;
	wire phi_n24_out1_ready;
	wire phi_n24_out1_valid;

	wire fork_20_clk;
	wire fork_20_rst;
	wire [31 : 0]fork_20_in1_data;
	wire fork_20_in1_ready;
	wire fork_20_in1_valid;
	wire [31 : 0]fork_20_out1_data;
	wire fork_20_out1_ready;
	wire fork_20_out1_valid;
	wire [31 : 0]fork_20_out2_data;
	wire fork_20_out2_ready;
	wire fork_20_out2_valid;

	wire fork_21_clk;
	wire fork_21_rst;
	wire [31 : 0]fork_21_in1_data;
	wire fork_21_in1_ready;
	wire fork_21_in1_valid;
	wire [31 : 0]fork_21_out1_data;
	wire fork_21_out1_ready;
	wire fork_21_out1_valid;
	wire [31 : 0]fork_21_out2_data;
	wire fork_21_out2_ready;
	wire fork_21_out2_valid;

	wire branch_27_clk;
	wire branch_27_rst;
	wire [31 : 0]branch_27_in1_data;
	wire branch_27_in1_ready;
	wire branch_27_in1_valid;
	wire [0 : 0]branch_27_in2_data;
	wire branch_27_in2_ready;
	wire branch_27_in2_valid;
	wire [31 : 0]branch_27_out1_data;
	wire branch_27_out1_ready;
	wire branch_27_out1_valid;
	wire [31 : 0]branch_27_out2_data;
	wire branch_27_out2_ready;
	wire branch_27_out2_valid;

	wire branch_28_clk;
	wire branch_28_rst;
	wire [31 : 0]branch_28_in1_data;
	wire branch_28_in1_ready;
	wire branch_28_in1_valid;
	wire [0 : 0]branch_28_in2_data;
	wire branch_28_in2_ready;
	wire branch_28_in2_valid;
	wire [31 : 0]branch_28_out1_data;
	wire branch_28_out1_ready;
	wire branch_28_out1_valid;
	wire [31 : 0]branch_28_out2_data;
	wire branch_28_out2_ready;
	wire branch_28_out2_valid;

	wire branch_29_clk;
	wire branch_29_rst;
	wire [31 : 0]branch_29_in1_data;
	wire branch_29_in1_ready;
	wire branch_29_in1_valid;
	wire [0 : 0]branch_29_in2_data;
	wire branch_29_in2_ready;
	wire branch_29_in2_valid;
	wire [31 : 0]branch_29_out1_data;
	wire branch_29_out1_ready;
	wire branch_29_out1_valid;
	wire [31 : 0]branch_29_out2_data;
	wire branch_29_out2_ready;
	wire branch_29_out2_valid;

	wire branch_30_clk;
	wire branch_30_rst;
	wire [9 : 0]branch_30_in1_data;
	wire branch_30_in1_ready;
	wire branch_30_in1_valid;
	wire [0 : 0]branch_30_in2_data;
	wire branch_30_in2_ready;
	wire branch_30_in2_valid;
	wire [9 : 0]branch_30_out1_data;
	wire branch_30_out1_ready;
	wire branch_30_out1_valid;
	wire [9 : 0]branch_30_out2_data;
	wire branch_30_out2_ready;
	wire branch_30_out2_valid;

	wire fork_36_clk;
	wire fork_36_rst;
	wire [0 : 0]fork_36_in1_data;
	wire fork_36_in1_ready;
	wire fork_36_in1_valid;
	wire [0 : 0]fork_36_out1_data;
	wire fork_36_out1_ready;
	wire fork_36_out1_valid;
	wire [0 : 0]fork_36_out2_data;
	wire fork_36_out2_ready;
	wire fork_36_out2_valid;
	wire [0 : 0]fork_36_out3_data;
	wire fork_36_out3_ready;
	wire fork_36_out3_valid;
	wire [0 : 0]fork_36_out4_data;
	wire fork_36_out4_ready;
	wire fork_36_out4_valid;
	wire [0 : 0]fork_36_out5_data;
	wire fork_36_out5_ready;
	wire fork_36_out5_valid;

	wire phiC_38_clk;
	wire phiC_38_rst;
	wire [0 : 0]phiC_38_in1_data;
	wire phiC_38_in1_ready;
	wire phiC_38_in1_valid;
	wire [0 : 0]phiC_38_out1_data;
	wire phiC_38_out1_ready;
	wire phiC_38_out1_valid;

	wire branchC_53_clk;
	wire branchC_53_rst;
	wire [0 : 0]branchC_53_in1_data;
	wire branchC_53_in1_ready;
	wire branchC_53_in1_valid;
	wire [0 : 0]branchC_53_in2_data;
	wire branchC_53_in2_ready;
	wire branchC_53_in2_valid;
	wire [0 : 0]branchC_53_out1_data;
	wire branchC_53_out1_ready;
	wire branchC_53_out1_valid;
	wire [0 : 0]branchC_53_out2_data;
	wire branchC_53_out2_ready;
	wire branchC_53_out2_valid;

	wire MC_kmpNext_clk;
	wire MC_kmpNext_rst;
	wire [31 : 0]MC_kmpNext_in1_data;
	wire MC_kmpNext_in1_ready;
	wire MC_kmpNext_in1_valid;
	wire [31 : 0]MC_kmpNext_in2_data;
	wire MC_kmpNext_in2_ready;
	wire MC_kmpNext_in2_valid;
	wire [31 : 0]MC_kmpNext_in3_data;
	wire MC_kmpNext_in3_ready;
	wire MC_kmpNext_in3_valid;
	wire [31 : 0]MC_kmpNext_in4_data;
	wire MC_kmpNext_in4_ready;
	wire MC_kmpNext_in4_valid;
	wire [31 : 0]MC_kmpNext_in5_data;
	wire MC_kmpNext_in5_ready;
	wire MC_kmpNext_in5_valid;
	wire [31 : 0]MC_kmpNext_in6_data;
	wire MC_kmpNext_in6_ready;
	wire MC_kmpNext_in6_valid;
	wire [31 : 0]MC_kmpNext_in7_data;
	wire MC_kmpNext_in7_ready;
	wire MC_kmpNext_in7_valid;
	wire [31 : 0]MC_kmpNext_in8_data;
	wire MC_kmpNext_in8_ready;
	wire MC_kmpNext_in8_valid;
	wire [31 : 0]MC_kmpNext_in9_data;
	wire MC_kmpNext_in9_ready;
	wire MC_kmpNext_in9_valid;
	wire [31 : 0]MC_kmpNext_out1_data;
	wire MC_kmpNext_out1_ready;
	wire MC_kmpNext_out1_valid;
	wire [31 : 0]MC_kmpNext_out2_data;
	wire MC_kmpNext_out2_ready;
	wire MC_kmpNext_out2_valid;
	wire [31 : 0]MC_kmpNext_out3_data;
	wire MC_kmpNext_out3_ready;
	wire MC_kmpNext_out3_valid;
	wire [0 : 0]MC_kmpNext_out4_data;
	wire MC_kmpNext_out4_ready;
	wire MC_kmpNext_out4_valid;

	wire MC_pattern_clk;
	wire MC_pattern_rst;
	wire [31 : 0]MC_pattern_in1_data;
	wire MC_pattern_in1_ready;
	wire MC_pattern_in1_valid;
	wire [31 : 0]MC_pattern_in2_data;
	wire MC_pattern_in2_ready;
	wire MC_pattern_in2_valid;
	wire [31 : 0]MC_pattern_in3_data;
	wire MC_pattern_in3_ready;
	wire MC_pattern_in3_valid;
	wire [31 : 0]MC_pattern_in4_data;
	wire MC_pattern_in4_ready;
	wire MC_pattern_in4_valid;
	wire [31 : 0]MC_pattern_in5_data;
	wire MC_pattern_in5_ready;
	wire MC_pattern_in5_valid;
	wire [31 : 0]MC_pattern_in6_data;
	wire MC_pattern_in6_ready;
	wire MC_pattern_in6_valid;
	wire [31 : 0]MC_pattern_in7_data;
	wire MC_pattern_in7_ready;
	wire MC_pattern_in7_valid;
	wire [31 : 0]MC_pattern_in8_data;
	wire MC_pattern_in8_ready;
	wire MC_pattern_in8_valid;
	wire [31 : 0]MC_pattern_out1_data;
	wire MC_pattern_out1_ready;
	wire MC_pattern_out1_valid;
	wire [31 : 0]MC_pattern_out2_data;
	wire MC_pattern_out2_ready;
	wire MC_pattern_out2_valid;
	wire [31 : 0]MC_pattern_out3_data;
	wire MC_pattern_out3_ready;
	wire MC_pattern_out3_valid;
	wire [31 : 0]MC_pattern_out4_data;
	wire MC_pattern_out4_ready;
	wire MC_pattern_out4_valid;
	wire [31 : 0]MC_pattern_out5_data;
	wire MC_pattern_out5_ready;
	wire MC_pattern_out5_valid;
	wire [0 : 0]MC_pattern_out6_data;
	wire MC_pattern_out6_ready;
	wire MC_pattern_out6_valid;

	wire MC_input_clk;
	wire MC_input_rst;
	wire [9 : 0]MC_input_in1_data;
	wire MC_input_in1_ready;
	wire MC_input_in1_valid;
	wire [31 : 0]MC_input_in2_data;
	wire MC_input_in2_ready;
	wire MC_input_in2_valid;
	wire [9 : 0]MC_input_in3_data;
	wire MC_input_in3_ready;
	wire MC_input_in3_valid;
	wire [31 : 0]MC_input_in4_data;
	wire MC_input_in4_ready;
	wire MC_input_in4_valid;
	wire [31 : 0]MC_input_out1_data;
	wire MC_input_out1_ready;
	wire MC_input_out1_valid;
	wire [0 : 0]MC_input_out2_data;
	wire MC_input_out2_ready;
	wire MC_input_out2_valid;

	wire sink_1_clk;
	wire sink_1_rst;
	wire [0 : 0]sink_1_in1_data;
	wire sink_1_in1_ready;
	wire sink_1_in1_valid;

	wire sink_2_clk;
	wire sink_2_rst;
	wire [0 : 0]sink_2_in1_data;
	wire sink_2_in1_ready;
	wire sink_2_in1_valid;

	wire sink_3_clk;
	wire sink_3_rst;
	wire [31 : 0]sink_3_in1_data;
	wire sink_3_in1_ready;
	wire sink_3_in1_valid;

	wire sink_4_clk;
	wire sink_4_rst;
	wire [31 : 0]sink_4_in1_data;
	wire sink_4_in1_ready;
	wire sink_4_in1_valid;

	wire sink_5_clk;
	wire sink_5_rst;
	wire [2 : 0]sink_5_in1_data;
	wire sink_5_in1_ready;
	wire sink_5_in1_valid;

	wire sink_6_clk;
	wire sink_6_rst;
	wire [31 : 0]sink_6_in1_data;
	wire sink_6_in1_ready;
	wire sink_6_in1_valid;

	wire sink_7_clk;
	wire sink_7_rst;
	wire [31 : 0]sink_7_in1_data;
	wire sink_7_in1_ready;
	wire sink_7_in1_valid;

	wire sink_8_clk;
	wire sink_8_rst;
	wire [31 : 0]sink_8_in1_data;
	wire sink_8_in1_ready;
	wire sink_8_in1_valid;

	wire sink_9_clk;
	wire sink_9_rst;
	wire [2 : 0]sink_9_in1_data;
	wire sink_9_in1_ready;
	wire sink_9_in1_valid;

	wire sink_10_clk;
	wire sink_10_rst;
	wire [31 : 0]sink_10_in1_data;
	wire sink_10_in1_ready;
	wire sink_10_in1_valid;

	wire sink_11_clk;
	wire sink_11_rst;
	wire [2 : 0]sink_11_in1_data;
	wire sink_11_in1_ready;
	wire sink_11_in1_valid;

	wire sink_12_clk;
	wire sink_12_rst;
	wire [0 : 0]sink_12_in1_data;
	wire sink_12_in1_ready;
	wire sink_12_in1_valid;

	wire sink_13_clk;
	wire sink_13_rst;
	wire [0 : 0]sink_13_in1_data;
	wire sink_13_in1_ready;
	wire sink_13_in1_valid;

	wire sink_14_clk;
	wire sink_14_rst;
	wire [0 : 0]sink_14_in1_data;
	wire sink_14_in1_ready;
	wire sink_14_in1_valid;

	wire sink_15_clk;
	wire sink_15_rst;
	wire [31 : 0]sink_15_in1_data;
	wire sink_15_in1_ready;
	wire sink_15_in1_valid;

	wire sink_16_clk;
	wire sink_16_rst;
	wire [31 : 0]sink_16_in1_data;
	wire sink_16_in1_ready;
	wire sink_16_in1_valid;

	wire sink_17_clk;
	wire sink_17_rst;
	wire [31 : 0]sink_17_in1_data;
	wire sink_17_in1_ready;
	wire sink_17_in1_valid;

	wire sink_18_clk;
	wire sink_18_rst;
	wire [9 : 0]sink_18_in1_data;
	wire sink_18_in1_ready;
	wire sink_18_in1_valid;

	wire sink_19_clk;
	wire sink_19_rst;
	wire [31 : 0]sink_19_in1_data;
	wire sink_19_in1_ready;
	wire sink_19_in1_valid;

	wire sink_20_clk;
	wire sink_20_rst;
	wire [31 : 0]sink_20_in1_data;
	wire sink_20_in1_ready;
	wire sink_20_in1_valid;

	wire sink_21_clk;
	wire sink_21_rst;
	wire [31 : 0]sink_21_in1_data;
	wire sink_21_in1_ready;
	wire sink_21_in1_valid;

	wire sink_22_clk;
	wire sink_22_rst;
	wire [9 : 0]sink_22_in1_data;
	wire sink_22_in1_ready;
	wire sink_22_in1_valid;

	wire sink_23_clk;
	wire sink_23_rst;
	wire [31 : 0]sink_23_in1_data;
	wire sink_23_in1_ready;
	wire sink_23_in1_valid;

	wire sink_24_clk;
	wire sink_24_rst;
	wire [31 : 0]sink_24_in1_data;
	wire sink_24_in1_ready;
	wire sink_24_in1_valid;

	wire sink_25_clk;
	wire sink_25_rst;
	wire [9 : 0]sink_25_in1_data;
	wire sink_25_in1_ready;
	wire sink_25_in1_valid;

	wire sink_26_clk;
	wire sink_26_rst;
	wire [31 : 0]sink_26_in1_data;
	wire sink_26_in1_ready;
	wire sink_26_in1_valid;

	wire sink_27_clk;
	wire sink_27_rst;
	wire [9 : 0]sink_27_in1_data;
	wire sink_27_in1_ready;
	wire sink_27_in1_valid;

	wire sink_28_clk;
	wire sink_28_rst;
	wire [0 : 0]sink_28_in1_data;
	wire sink_28_in1_ready;
	wire sink_28_in1_valid;

	wire sink_29_clk;
	wire sink_29_rst;
	wire [0 : 0]sink_29_in1_data;
	wire sink_29_in1_ready;
	wire sink_29_in1_valid;

	wire sink_30_clk;
	wire sink_30_rst;
	wire [0 : 0]sink_30_in1_data;
	wire sink_30_in1_ready;
	wire sink_30_in1_valid;

	wire sink_31_clk;
	wire sink_31_rst;
	wire [0 : 0]sink_31_in1_data;
	wire sink_31_in1_ready;
	wire sink_31_in1_valid;

	wire sink_32_clk;
	wire sink_32_rst;
	wire [0 : 0]sink_32_in1_data;
	wire sink_32_in1_ready;
	wire sink_32_in1_valid;

	wire sink_33_clk;
	wire sink_33_rst;
	wire [0 : 0]sink_33_in1_data;
	wire sink_33_in1_ready;
	wire sink_33_in1_valid;

	wire sink_34_clk;
	wire sink_34_rst;
	wire [0 : 0]sink_34_in1_data;
	wire sink_34_in1_ready;
	wire sink_34_in1_valid;

	wire Buffer_100_clk;
	wire Buffer_100_rst;
	wire [31 : 0]Buffer_100_in1_data;
	wire Buffer_100_in1_ready;
	wire Buffer_100_in1_valid;
	wire [31 : 0]Buffer_100_out1_data;
	wire Buffer_100_out1_ready;
	wire Buffer_100_out1_valid;

	wire Buffer_101_clk;
	wire Buffer_101_rst;
	wire [31 : 0]Buffer_101_in1_data;
	wire Buffer_101_in1_ready;
	wire Buffer_101_in1_valid;
	wire [31 : 0]Buffer_101_out1_data;
	wire Buffer_101_out1_ready;
	wire Buffer_101_out1_valid;

	wire Buffer_102_clk;
	wire Buffer_102_rst;
	wire [31 : 0]Buffer_102_in1_data;
	wire Buffer_102_in1_ready;
	wire Buffer_102_in1_valid;
	wire [31 : 0]Buffer_102_out1_data;
	wire Buffer_102_out1_ready;
	wire Buffer_102_out1_valid;

	wire Buffer_103_clk;
	wire Buffer_103_rst;
	wire [31 : 0]Buffer_103_in1_data;
	wire Buffer_103_in1_ready;
	wire Buffer_103_in1_valid;
	wire [31 : 0]Buffer_103_out1_data;
	wire Buffer_103_out1_ready;
	wire Buffer_103_out1_valid;

	wire Buffer_104_clk;
	wire Buffer_104_rst;
	wire [31 : 0]Buffer_104_in1_data;
	wire Buffer_104_in1_ready;
	wire Buffer_104_in1_valid;
	wire [31 : 0]Buffer_104_out1_data;
	wire Buffer_104_out1_ready;
	wire Buffer_104_out1_valid;

	wire Buffer_105_clk;
	wire Buffer_105_rst;
	wire [31 : 0]Buffer_105_in1_data;
	wire Buffer_105_in1_ready;
	wire Buffer_105_in1_valid;
	wire [31 : 0]Buffer_105_out1_data;
	wire Buffer_105_out1_ready;
	wire Buffer_105_out1_valid;

	wire Buffer_106_clk;
	wire Buffer_106_rst;
	wire [31 : 0]Buffer_106_in1_data;
	wire Buffer_106_in1_ready;
	wire Buffer_106_in1_valid;
	wire [31 : 0]Buffer_106_out1_data;
	wire Buffer_106_out1_ready;
	wire Buffer_106_out1_valid;

	wire Buffer_107_clk;
	wire Buffer_107_rst;
	wire [31 : 0]Buffer_107_in1_data;
	wire Buffer_107_in1_ready;
	wire Buffer_107_in1_valid;
	wire [31 : 0]Buffer_107_out1_data;
	wire Buffer_107_out1_ready;
	wire Buffer_107_out1_valid;

	wire Buffer_108_clk;
	wire Buffer_108_rst;
	wire [31 : 0]Buffer_108_in1_data;
	wire Buffer_108_in1_ready;
	wire Buffer_108_in1_valid;
	wire [31 : 0]Buffer_108_out1_data;
	wire Buffer_108_out1_ready;
	wire Buffer_108_out1_valid;

	wire Buffer_109_clk;
	wire Buffer_109_rst;
	wire [31 : 0]Buffer_109_in1_data;
	wire Buffer_109_in1_ready;
	wire Buffer_109_in1_valid;
	wire [31 : 0]Buffer_109_out1_data;
	wire Buffer_109_out1_ready;
	wire Buffer_109_out1_valid;

	wire Buffer_110_clk;
	wire Buffer_110_rst;
	wire [31 : 0]Buffer_110_in1_data;
	wire Buffer_110_in1_ready;
	wire Buffer_110_in1_valid;
	wire [31 : 0]Buffer_110_out1_data;
	wire Buffer_110_out1_ready;
	wire Buffer_110_out1_valid;

	wire Buffer_111_clk;
	wire Buffer_111_rst;
	wire [31 : 0]Buffer_111_in1_data;
	wire Buffer_111_in1_ready;
	wire Buffer_111_in1_valid;
	wire [31 : 0]Buffer_111_out1_data;
	wire Buffer_111_out1_ready;
	wire Buffer_111_out1_valid;

	wire Buffer_112_clk;
	wire Buffer_112_rst;
	wire [31 : 0]Buffer_112_in1_data;
	wire Buffer_112_in1_ready;
	wire Buffer_112_in1_valid;
	wire [31 : 0]Buffer_112_out1_data;
	wire Buffer_112_out1_ready;
	wire Buffer_112_out1_valid;

	wire Buffer_113_clk;
	wire Buffer_113_rst;
	wire [31 : 0]Buffer_113_in1_data;
	wire Buffer_113_in1_ready;
	wire Buffer_113_in1_valid;
	wire [31 : 0]Buffer_113_out1_data;
	wire Buffer_113_out1_ready;
	wire Buffer_113_out1_valid;

	wire Buffer_114_clk;
	wire Buffer_114_rst;
	wire [31 : 0]Buffer_114_in1_data;
	wire Buffer_114_in1_ready;
	wire Buffer_114_in1_valid;
	wire [31 : 0]Buffer_114_out1_data;
	wire Buffer_114_out1_ready;
	wire Buffer_114_out1_valid;

	wire Buffer_115_clk;
	wire Buffer_115_rst;
	wire [31 : 0]Buffer_115_in1_data;
	wire Buffer_115_in1_ready;
	wire Buffer_115_in1_valid;
	wire [31 : 0]Buffer_115_out1_data;
	wire Buffer_115_out1_ready;
	wire Buffer_115_out1_valid;



	assign phi_1_clk = clk;
	assign phi_1_rst = rst;
	assign branch_2_in1_data = phi_1_out1_data;
	assign branch_2_in1_valid = phi_1_out1_valid;
	assign phi_1_out1_ready = branch_2_in1_ready;

	assign phi_2_clk = clk;
	assign phi_2_rst = rst;
	assign fork_0_in1_data = phi_2_out1_data;
	assign fork_0_in1_valid = phi_2_out1_valid;
	assign phi_2_out1_ready = fork_0_in1_ready;

	assign load_5_clk = clk;
	assign load_5_rst = rst;
	assign branch_3_in1_data = load_5_out1_data;
	assign branch_3_in1_valid = load_5_out1_valid;
	assign load_5_out1_ready = branch_3_in1_ready;
	assign MC_pattern_in1_data = load_5_out2_data;
	assign MC_pattern_in1_valid = load_5_out2_valid;
	assign load_5_out2_ready = MC_pattern_in1_ready;

	assign brCst_block2_clk = clk;
	assign brCst_block2_rst = rst;
	assign fork_28_in1_data = brCst_block2_out1_data;
	assign fork_28_in1_valid = brCst_block2_out1_valid;
	assign brCst_block2_out1_ready = fork_28_in1_ready;

	assign fork_0_clk = clk;
	assign fork_0_rst = rst;
	assign load_5_in2_data = fork_0_out1_data;
	assign load_5_in2_valid = fork_0_out1_valid;
	assign fork_0_out1_ready = load_5_in2_ready;
	assign branch_4_in1_data = fork_0_out2_data;
	assign branch_4_in1_valid = fork_0_out2_valid;
	assign fork_0_out2_ready = branch_4_in1_ready;

	assign branch_2_clk = clk;
	assign branch_2_rst = rst;
	assign phi_7_in2_data = branch_2_out1_data;
	assign phi_7_in2_valid = branch_2_out1_valid;
	assign branch_2_out1_ready = phi_7_in2_ready;
	assign sink_3_in1_data = branch_2_out2_data;
	assign sink_3_in1_valid = branch_2_out2_valid;
	assign branch_2_out2_ready = sink_3_in1_ready;

	assign branch_3_clk = clk;
	assign branch_3_rst = rst;
	assign phi_n6_in1_data = branch_3_out1_data;
	assign phi_n6_in1_valid = branch_3_out1_valid;
	assign branch_3_out1_ready = phi_n6_in1_ready;
	assign sink_4_in1_data = branch_3_out2_data;
	assign sink_4_in1_valid = branch_3_out2_valid;
	assign branch_3_out2_ready = sink_4_in1_ready;

	assign branch_4_clk = clk;
	assign branch_4_rst = rst;
	assign phi_n7_in1_data = branch_4_out1_data;
	assign phi_n7_in1_valid = branch_4_out1_valid;
	assign branch_4_out1_ready = phi_n7_in1_ready;
	assign sink_5_in1_data = branch_4_out2_data;
	assign sink_5_in1_valid = branch_4_out2_valid;
	assign branch_4_out2_ready = sink_5_in1_ready;

	assign fork_28_clk = clk;
	assign fork_28_rst = rst;
	assign branch_4_in2_data = fork_28_out1_data;
	assign branch_4_in2_valid = fork_28_out1_valid;
	assign fork_28_out1_ready = branch_4_in2_ready;
	assign branch_3_in2_data = fork_28_out2_data;
	assign branch_3_in2_valid = fork_28_out2_valid;
	assign fork_28_out2_ready = branch_3_in2_ready;
	assign branch_2_in2_data = fork_28_out3_data;
	assign branch_2_in2_valid = fork_28_out3_valid;
	assign fork_28_out3_ready = branch_2_in2_ready;
	assign branchC_45_in2_data = fork_28_out4_data;
	assign branchC_45_in2_valid = fork_28_out4_valid;
	assign fork_28_out4_ready = branchC_45_in2_ready;

	assign phiC_30_clk = clk;
	assign phiC_30_rst = rst;
	assign forkC_43_in1_data = phiC_30_out1_data;
	assign forkC_43_in1_valid = phiC_30_out1_valid;
	assign phiC_30_out1_ready = forkC_43_in1_ready;
	assign fork_57_in1_data = phiC_30_out2_data;
	assign fork_57_in1_valid = phiC_30_out2_valid;
	assign phiC_30_out2_ready = fork_57_in1_ready;

	assign forkC_43_clk = clk;
	assign forkC_43_rst = rst;
	assign branchC_45_in1_data = forkC_43_out1_data;
	assign branchC_45_in1_valid = forkC_43_out1_valid;
	assign forkC_43_out1_ready = branchC_45_in1_ready;
	assign brCst_block2_in1_data = forkC_43_out2_data;
	assign brCst_block2_in1_valid = forkC_43_out2_valid;
	assign forkC_43_out2_ready = brCst_block2_in1_ready;

	assign branchC_45_clk = clk;
	assign branchC_45_rst = rst;
	assign phiC_31_in1_data = branchC_45_out1_data;
	assign phiC_31_in1_valid = branchC_45_out1_valid;
	assign branchC_45_out1_ready = phiC_31_in1_ready;
	assign sink_29_in1_data = branchC_45_out2_data;
	assign sink_29_in1_valid = branchC_45_out2_valid;
	assign branchC_45_out2_ready = sink_29_in1_ready;

	assign fork_57_clk = clk;
	assign fork_57_rst = rst;
	assign phi_1_in1_data = fork_57_out1_data;
	assign phi_1_in1_valid = fork_57_out1_valid;
	assign fork_57_out1_ready = phi_1_in1_ready;
	assign phi_2_in1_data = fork_57_out2_data;
	assign phi_2_in1_valid = fork_57_out2_valid;
	assign fork_57_out2_ready = phi_2_in1_ready;

	assign phi_31_clk = clk;
	assign phi_31_rst = rst;
	assign branch_21_in1_data = phi_31_out1_data;
	assign branch_21_in1_valid = phi_31_out1_valid;
	assign phi_31_out1_ready = branch_21_in1_ready;

	assign phi_32_clk = clk;
	assign phi_32_rst = rst;
	assign branch_19_in1_data = phi_32_out1_data;
	assign branch_19_in1_valid = phi_32_out1_valid;
	assign phi_32_out1_ready = branch_19_in1_ready;

	assign phi_33_clk = clk;
	assign phi_33_rst = rst;
	assign fork_4_in1_data = phi_33_out1_data;
	assign fork_4_in1_valid = phi_33_out1_valid;
	assign phi_33_out1_ready = fork_4_in1_ready;

	assign load_36_clk = clk;
	assign load_36_rst = rst;
	assign branch_20_in1_data = load_36_out1_data;
	assign branch_20_in1_valid = load_36_out1_valid;
	assign load_36_out1_ready = branch_20_in1_ready;
	assign MC_input_in1_data = load_36_out2_data;
	assign MC_input_in1_valid = load_36_out2_valid;
	assign load_36_out2_ready = MC_input_in1_ready;

	assign brCst_block8_clk = clk;
	assign brCst_block8_rst = rst;
	assign fork_34_in1_data = brCst_block8_out1_data;
	assign fork_34_in1_valid = brCst_block8_out1_valid;
	assign brCst_block8_out1_ready = fork_34_in1_ready;

	assign fork_4_clk = clk;
	assign fork_4_rst = rst;
	assign load_36_in2_data = fork_4_out1_data;
	assign load_36_in2_valid = fork_4_out1_valid;
	assign fork_4_out1_ready = load_36_in2_ready;
	assign branch_22_in1_data = fork_4_out2_data;
	assign branch_22_in1_valid = fork_4_out2_valid;
	assign fork_4_out2_ready = branch_22_in1_ready;

	assign branch_19_clk = clk;
	assign branch_19_rst = rst;
	assign phi_38_in2_data = branch_19_out1_data;
	assign phi_38_in2_valid = branch_19_out1_valid;
	assign branch_19_out1_ready = phi_38_in2_ready;
	assign sink_15_in1_data = branch_19_out2_data;
	assign sink_15_in1_valid = branch_19_out2_valid;
	assign branch_19_out2_ready = sink_15_in1_ready;

	assign branch_20_clk = clk;
	assign branch_20_rst = rst;
	assign phi_n10_in1_data = branch_20_out1_data;
	assign phi_n10_in1_valid = branch_20_out1_valid;
	assign branch_20_out1_ready = phi_n10_in1_ready;
	assign sink_16_in1_data = branch_20_out2_data;
	assign sink_16_in1_valid = branch_20_out2_valid;
	assign branch_20_out2_ready = sink_16_in1_ready;

	assign branch_21_clk = clk;
	assign branch_21_rst = rst;
	assign phi_n11_in1_data = branch_21_out1_data;
	assign phi_n11_in1_valid = branch_21_out1_valid;
	assign branch_21_out1_ready = phi_n11_in1_ready;
	assign sink_17_in1_data = branch_21_out2_data;
	assign sink_17_in1_valid = branch_21_out2_valid;
	assign branch_21_out2_ready = sink_17_in1_ready;

	assign branch_22_clk = clk;
	assign branch_22_rst = rst;
	assign phi_n12_in1_data = branch_22_out1_data;
	assign phi_n12_in1_valid = branch_22_out1_valid;
	assign branch_22_out1_ready = phi_n12_in1_ready;
	assign sink_18_in1_data = branch_22_out2_data;
	assign sink_18_in1_valid = branch_22_out2_valid;
	assign branch_22_out2_ready = sink_18_in1_ready;

	assign fork_34_clk = clk;
	assign fork_34_rst = rst;
	assign branch_22_in2_data = fork_34_out1_data;
	assign branch_22_in2_valid = fork_34_out1_valid;
	assign fork_34_out1_ready = branch_22_in2_ready;
	assign branch_21_in2_data = fork_34_out2_data;
	assign branch_21_in2_valid = fork_34_out2_valid;
	assign fork_34_out2_ready = branch_21_in2_ready;
	assign branch_20_in2_data = fork_34_out3_data;
	assign branch_20_in2_valid = fork_34_out3_valid;
	assign fork_34_out3_ready = branch_20_in2_ready;
	assign branch_19_in2_data = fork_34_out4_data;
	assign branch_19_in2_valid = fork_34_out4_valid;
	assign fork_34_out4_ready = branch_19_in2_ready;
	assign branchC_51_in2_data = fork_34_out5_data;
	assign branchC_51_in2_valid = fork_34_out5_valid;
	assign fork_34_out5_ready = branchC_51_in2_ready;

	assign phiC_36_clk = clk;
	assign phiC_36_rst = rst;
	assign forkC_49_in1_data = phiC_36_out1_data;
	assign forkC_49_in1_valid = phiC_36_out1_valid;
	assign phiC_36_out1_ready = forkC_49_in1_ready;
	assign fork_59_in1_data = phiC_36_out2_data;
	assign fork_59_in1_valid = phiC_36_out2_valid;
	assign phiC_36_out2_ready = fork_59_in1_ready;

	assign forkC_49_clk = clk;
	assign forkC_49_rst = rst;
	assign branchC_51_in1_data = forkC_49_out1_data;
	assign branchC_51_in1_valid = forkC_49_out1_valid;
	assign forkC_49_out1_ready = branchC_51_in1_ready;
	assign brCst_block8_in1_data = forkC_49_out2_data;
	assign brCst_block8_in1_valid = forkC_49_out2_valid;
	assign forkC_49_out2_ready = brCst_block8_in1_ready;

	assign branchC_51_clk = clk;
	assign branchC_51_rst = rst;
	assign phiC_37_in1_data = branchC_51_out1_data;
	assign phiC_37_in1_valid = branchC_51_out1_valid;
	assign branchC_51_out1_ready = phiC_37_in1_ready;
	assign sink_32_in1_data = branchC_51_out2_data;
	assign sink_32_in1_valid = branchC_51_out2_valid;
	assign branchC_51_out2_ready = sink_32_in1_ready;

	assign fork_59_clk = clk;
	assign fork_59_rst = rst;
	assign phi_31_in1_data = fork_59_out1_data;
	assign phi_31_in1_valid = fork_59_out1_valid;
	assign fork_59_out1_ready = phi_31_in1_ready;
	assign phi_32_in1_data = fork_59_out2_data;
	assign phi_32_in1_valid = fork_59_out2_valid;
	assign fork_59_out2_ready = phi_32_in1_ready;
	assign phi_33_in1_data = fork_59_out3_data;
	assign phi_33_in1_valid = fork_59_out3_valid;
	assign fork_59_out3_ready = phi_33_in1_ready;

	assign load_48_clk = clk;
	assign load_48_rst = rst;
	assign branch_31_in1_data = load_48_out1_data;
	assign branch_31_in1_valid = load_48_out1_valid;
	assign load_48_out1_ready = branch_31_in1_ready;
	assign MC_kmpNext_in8_data = load_48_out2_data;
	assign MC_kmpNext_in8_valid = load_48_out2_valid;
	assign load_48_out2_ready = MC_kmpNext_in8_ready;

	assign brCst_block11_clk = clk;
	assign brCst_block11_rst = rst;
	assign fork_37_in1_data = brCst_block11_out1_data;
	assign fork_37_in1_valid = brCst_block11_out1_valid;
	assign brCst_block11_out1_ready = fork_37_in1_ready;

	assign phi_n17_clk = clk;
	assign phi_n17_rst = rst;
	assign load_48_in2_data = phi_n17_out1_data;
	assign load_48_in2_valid = phi_n17_out1_valid;
	assign phi_n17_out1_ready = load_48_in2_ready;

	assign phi_n18_clk = clk;
	assign phi_n18_rst = rst;
	assign branch_32_in1_data = phi_n18_out1_data;
	assign branch_32_in1_valid = phi_n18_out1_valid;
	assign phi_n18_out1_ready = branch_32_in1_ready;

	assign phi_n19_clk = clk;
	assign phi_n19_rst = rst;
	assign branch_33_in1_data = phi_n19_out1_data;
	assign branch_33_in1_valid = phi_n19_out1_valid;
	assign phi_n19_out1_ready = branch_33_in1_ready;

	assign phi_n20_clk = clk;
	assign phi_n20_rst = rst;
	assign branch_34_in1_data = phi_n20_out1_data;
	assign branch_34_in1_valid = phi_n20_out1_valid;
	assign phi_n20_out1_ready = branch_34_in1_ready;

	assign branch_31_clk = clk;
	assign branch_31_rst = rst;
	assign Buffer_107_in1_data = branch_31_out1_data;
	assign Buffer_107_in1_valid = branch_31_out1_valid;
	assign branch_31_out1_ready = Buffer_107_in1_ready;
	assign sink_19_in1_data = branch_31_out2_data;
	assign sink_19_in1_valid = branch_31_out2_valid;
	assign branch_31_out2_ready = sink_19_in1_ready;

	assign branch_32_clk = clk;
	assign branch_32_rst = rst;
	assign Buffer_108_in1_data = branch_32_out1_data;
	assign Buffer_108_in1_valid = branch_32_out1_valid;
	assign branch_32_out1_ready = Buffer_108_in1_ready;
	assign sink_20_in1_data = branch_32_out2_data;
	assign sink_20_in1_valid = branch_32_out2_valid;
	assign branch_32_out2_ready = sink_20_in1_ready;

	assign branch_33_clk = clk;
	assign branch_33_rst = rst;
	assign Buffer_109_in1_data = branch_33_out1_data;
	assign Buffer_109_in1_valid = branch_33_out1_valid;
	assign branch_33_out1_ready = Buffer_109_in1_ready;
	assign sink_21_in1_data = branch_33_out2_data;
	assign sink_21_in1_valid = branch_33_out2_valid;
	assign branch_33_out2_ready = sink_21_in1_ready;

	assign branch_34_clk = clk;
	assign branch_34_rst = rst;
	assign Buffer_110_in1_data = branch_34_out1_data;
	assign Buffer_110_in1_valid = branch_34_out1_valid;
	assign branch_34_out1_ready = Buffer_110_in1_ready;
	assign sink_22_in1_data = branch_34_out2_data;
	assign sink_22_in1_valid = branch_34_out2_valid;
	assign branch_34_out2_ready = sink_22_in1_ready;

	assign fork_37_clk = clk;
	assign fork_37_rst = rst;
	assign branch_34_in2_data = fork_37_out1_data;
	assign branch_34_in2_valid = fork_37_out1_valid;
	assign fork_37_out1_ready = branch_34_in2_ready;
	assign branch_33_in2_data = fork_37_out2_data;
	assign branch_33_in2_valid = fork_37_out2_valid;
	assign fork_37_out2_ready = branch_33_in2_ready;
	assign branch_32_in2_data = fork_37_out3_data;
	assign branch_32_in2_valid = fork_37_out3_valid;
	assign fork_37_out3_ready = branch_32_in2_ready;
	assign branch_31_in2_data = fork_37_out4_data;
	assign branch_31_in2_valid = fork_37_out4_valid;
	assign fork_37_out4_ready = branch_31_in2_ready;
	assign branchC_54_in2_data = fork_37_out5_data;
	assign branchC_54_in2_valid = fork_37_out5_valid;
	assign fork_37_out5_ready = branchC_54_in2_ready;

	assign phiC_39_clk = clk;
	assign phiC_39_rst = rst;
	assign forkC_52_in1_data = phiC_39_out1_data;
	assign forkC_52_in1_valid = phiC_39_out1_valid;
	assign phiC_39_out1_ready = forkC_52_in1_ready;

	assign forkC_52_clk = clk;
	assign forkC_52_rst = rst;
	assign branchC_54_in1_data = forkC_52_out1_data;
	assign branchC_54_in1_valid = forkC_52_out1_valid;
	assign forkC_52_out1_ready = branchC_54_in1_ready;
	assign brCst_block11_in1_data = forkC_52_out2_data;
	assign brCst_block11_in1_valid = forkC_52_out2_valid;
	assign forkC_52_out2_ready = brCst_block11_in1_ready;

	assign branchC_54_clk = clk;
	assign branchC_54_rst = rst;
	assign Buffer_111_in1_data = branchC_54_out1_data;
	assign Buffer_111_in1_valid = branchC_54_out1_valid;
	assign branchC_54_out1_ready = Buffer_111_in1_ready;
	assign sink_33_in1_data = branchC_54_out2_data;
	assign sink_33_in1_valid = branchC_54_out2_valid;
	assign branchC_54_out2_ready = sink_33_in1_ready;

	assign load_52_clk = clk;
	assign load_52_rst = rst;
	assign icmp_53_in1_data = load_52_out1_data;
	assign icmp_53_in1_valid = load_52_out1_valid;
	assign load_52_out1_ready = icmp_53_in1_ready;
	assign MC_pattern_in5_data = load_52_out2_data;
	assign MC_pattern_in5_valid = load_52_out2_valid;
	assign load_52_out2_ready = MC_pattern_in5_ready;

	assign icmp_53_clk = clk;
	assign icmp_53_rst = rst;
	assign zext_54_in1_data = icmp_53_out1_data;
	assign zext_54_in1_valid = icmp_53_out1_valid;
	assign icmp_53_out1_ready = zext_54_in1_ready;

	assign zext_54_clk = clk;
	assign zext_54_rst = rst;
	assign add_55_in2_data = zext_54_out1_data;
	assign add_55_in2_valid = zext_54_out1_valid;
	assign zext_54_out1_ready = add_55_in2_ready;

	assign add_55_clk = clk;
	assign add_55_rst = rst;
	assign fork_6_in1_data = add_55_out1_data;
	assign fork_6_in1_valid = add_55_out1_valid;
	assign add_55_out1_ready = fork_6_in1_ready;

	assign cst_10_clk = clk;
	assign cst_10_rst = rst;
	assign icmp_56_in2_data = cst_10_out1_data;
	assign icmp_56_in2_valid = cst_10_out1_valid;
	assign cst_10_out1_ready = icmp_56_in2_ready;

	assign icmp_56_clk = clk;
	assign icmp_56_rst = rst;
	assign fork_38_in1_data = icmp_56_out1_data;
	assign fork_38_in1_valid = icmp_56_out1_valid;
	assign icmp_56_out1_ready = fork_38_in1_ready;

	assign phi_n25_clk = clk;
	assign phi_n25_rst = rst;
	assign fork_24_in1_data = phi_n25_out1_data;
	assign fork_24_in1_valid = phi_n25_out1_valid;
	assign phi_n25_out1_ready = fork_24_in1_ready;

	assign phi_n26_clk = clk;
	assign phi_n26_rst = rst;
	assign icmp_53_in2_data = phi_n26_out1_data;
	assign icmp_53_in2_valid = phi_n26_out1_valid;
	assign phi_n26_out1_ready = icmp_53_in2_ready;

	assign phi_n27_clk = clk;
	assign phi_n27_rst = rst;
	assign branch_36_in1_data = phi_n27_out1_data;
	assign branch_36_in1_valid = phi_n27_out1_valid;
	assign phi_n27_out1_ready = branch_36_in1_ready;

	assign phi_n28_clk = clk;
	assign phi_n28_rst = rst;
	assign branch_37_in1_data = phi_n28_out1_data;
	assign branch_37_in1_valid = phi_n28_out1_valid;
	assign phi_n28_out1_ready = branch_37_in1_ready;

	assign fork_6_clk = clk;
	assign fork_6_rst = rst;
	assign icmp_56_in1_data = fork_6_out1_data;
	assign icmp_56_in1_valid = fork_6_out1_valid;
	assign fork_6_out1_ready = icmp_56_in1_ready;
	assign branch_35_in1_data = fork_6_out2_data;
	assign branch_35_in1_valid = fork_6_out2_valid;
	assign fork_6_out2_ready = branch_35_in1_ready;

	assign fork_24_clk = clk;
	assign fork_24_rst = rst;
	assign load_52_in2_data = fork_24_out1_data;
	assign load_52_in2_valid = fork_24_out1_valid;
	assign fork_24_out1_ready = load_52_in2_ready;
	assign add_55_in1_data = fork_24_out2_data;
	assign add_55_in1_valid = fork_24_out2_valid;
	assign fork_24_out2_ready = add_55_in1_ready;

	assign branch_35_clk = clk;
	assign branch_35_rst = rst;
	assign phi_n14_in1_data = branch_35_out1_data;
	assign phi_n14_in1_valid = branch_35_out1_valid;
	assign branch_35_out1_ready = phi_n14_in1_ready;
	assign phi_64_in2_data = branch_35_out2_data;
	assign phi_64_in2_valid = branch_35_out2_valid;
	assign branch_35_out2_ready = phi_64_in2_ready;

	assign branch_36_clk = clk;
	assign branch_36_rst = rst;
	assign phi_n13_in1_data = branch_36_out1_data;
	assign phi_n13_in1_valid = branch_36_out1_valid;
	assign branch_36_out1_ready = phi_n13_in1_ready;
	assign phi_65_in2_data = branch_36_out2_data;
	assign phi_65_in2_valid = branch_36_out2_valid;
	assign branch_36_out2_ready = phi_65_in2_ready;

	assign branch_37_clk = clk;
	assign branch_37_rst = rst;
	assign phi_n15_in1_data = branch_37_out1_data;
	assign phi_n15_in1_valid = branch_37_out1_valid;
	assign branch_37_out1_ready = phi_n15_in1_ready;
	assign phi_n16_in1_data = branch_37_out2_data;
	assign phi_n16_in1_valid = branch_37_out2_valid;
	assign branch_37_out2_ready = phi_n16_in1_ready;

	assign fork_38_clk = clk;
	assign fork_38_rst = rst;
	assign branch_37_in2_data = fork_38_out1_data;
	assign branch_37_in2_valid = fork_38_out1_valid;
	assign fork_38_out1_ready = branch_37_in2_ready;
	assign branch_36_in2_data = fork_38_out2_data;
	assign branch_36_in2_valid = fork_38_out2_valid;
	assign fork_38_out2_ready = branch_36_in2_ready;
	assign branch_35_in2_data = fork_38_out3_data;
	assign branch_35_in2_valid = fork_38_out3_valid;
	assign fork_38_out3_ready = branch_35_in2_ready;
	assign branchC_55_in2_data = fork_38_out4_data;
	assign branchC_55_in2_valid = fork_38_out4_valid;
	assign fork_38_out4_ready = branchC_55_in2_ready;

	assign phiC_40_clk = clk;
	assign phiC_40_rst = rst;
	assign branchC_55_in1_data = phiC_40_out1_data;
	assign branchC_55_in1_valid = phiC_40_out1_valid;
	assign phiC_40_out1_ready = branchC_55_in1_ready;

	assign branchC_55_clk = clk;
	assign branchC_55_rst = rst;
	assign phiC_41_in1_data = branchC_55_out1_data;
	assign phiC_41_in1_valid = branchC_55_out1_valid;
	assign branchC_55_out1_ready = phiC_41_in1_ready;
	assign phiC_42_in1_data = branchC_55_out2_data;
	assign phiC_42_in1_valid = branchC_55_out2_valid;
	assign branchC_55_out2_ready = phiC_42_in1_ready;

	assign source_4_clk = clk;
	assign source_4_rst = rst;
	assign cst_10_in1_data = source_4_out1_data;
	assign cst_10_in1_valid = source_4_out1_valid;
	assign source_4_out1_ready = cst_10_in1_ready;

	assign cst_0_clk = clk;
	assign cst_0_rst = rst;
	assign store_0_in1_data = cst_0_out1_data;
	assign store_0_in1_valid = cst_0_out1_valid;
	assign cst_0_out1_ready = store_0_in1_ready;

	assign store_0_clk = clk;
	assign store_0_rst = rst;
	assign MC_kmpNext_in4_data = store_0_out1_data;
	assign MC_kmpNext_in4_valid = store_0_out1_valid;
	assign store_0_out1_ready = MC_kmpNext_in4_ready;
	assign MC_kmpNext_in3_data = store_0_out2_data;
	assign MC_kmpNext_in3_valid = store_0_out2_valid;
	assign store_0_out2_ready = MC_kmpNext_in3_ready;

	assign brCst_block1_clk = clk;
	assign brCst_block1_rst = rst;
	assign fork_27_in1_data = brCst_block1_out1_data;
	assign fork_27_in1_valid = brCst_block1_out1_valid;
	assign brCst_block1_out1_ready = fork_27_in1_ready;

	assign cst_1_clk = clk;
	assign cst_1_rst = rst;
	assign branch_0_in1_data = cst_1_out1_data;
	assign branch_0_in1_valid = cst_1_out1_valid;
	assign cst_1_out1_ready = branch_0_in1_ready;

	assign cst_2_clk = clk;
	assign cst_2_rst = rst;
	assign branch_1_in1_data = cst_2_out1_data;
	assign branch_1_in1_valid = cst_2_out1_valid;
	assign cst_2_out1_ready = branch_1_in1_ready;

	assign cst_15_clk = clk;
	assign cst_15_rst = rst;
	assign store_0_in2_data = cst_15_out1_data;
	assign store_0_in2_valid = cst_15_out1_valid;
	assign cst_15_out1_ready = store_0_in2_ready;

	assign branch_0_clk = clk;
	assign branch_0_rst = rst;
	assign phi_1_in2_data = branch_0_out1_data;
	assign phi_1_in2_valid = branch_0_out1_valid;
	assign branch_0_out1_ready = phi_1_in2_ready;
	assign sink_1_in1_data = branch_0_out2_data;
	assign sink_1_in1_valid = branch_0_out2_valid;
	assign branch_0_out2_ready = sink_1_in1_ready;

	assign branch_1_clk = clk;
	assign branch_1_rst = rst;
	assign phi_2_in2_data = branch_1_out1_data;
	assign phi_2_in2_valid = branch_1_out1_valid;
	assign branch_1_out1_ready = phi_2_in2_ready;
	assign sink_2_in1_data = branch_1_out2_data;
	assign sink_2_in1_valid = branch_1_out2_valid;
	assign branch_1_out2_ready = sink_2_in1_ready;

	assign fork_27_clk = clk;
	assign fork_27_rst = rst;
	assign branch_1_in2_data = fork_27_out1_data;
	assign branch_1_in2_valid = fork_27_out1_valid;
	assign fork_27_out1_ready = branch_1_in2_ready;
	assign branch_0_in2_data = fork_27_out2_data;
	assign branch_0_in2_valid = fork_27_out2_valid;
	assign fork_27_out2_ready = branch_0_in2_ready;
	assign branchC_44_in2_data = fork_27_out3_data;
	assign branchC_44_in2_valid = fork_27_out3_valid;
	assign fork_27_out3_ready = branchC_44_in2_ready;

	assign cst_16_clk = clk;
	assign cst_16_rst = rst;
	assign MC_kmpNext_in1_data = cst_16_out1_data;
	assign MC_kmpNext_in1_valid = cst_16_out1_valid;
	assign cst_16_out1_ready = MC_kmpNext_in1_ready;

	assign start_0_clk = clk;
	assign start_0_rst = rst;
	assign start_0_in1_data = start_in;
	assign start_0_in1_valid = start_valid;
	assign start_ready = start_0_in1_ready;
	assign forkC_42_in1_data = start_0_out1_data;
	assign forkC_42_in1_valid = start_0_out1_valid;
	assign start_0_out1_ready = forkC_42_in1_ready;

	assign forkC_42_clk = clk;
	assign forkC_42_rst = rst;
	assign cst_0_in1_data = forkC_42_out1_data;
	assign cst_0_in1_valid = forkC_42_out1_valid;
	assign forkC_42_out1_ready = cst_0_in1_ready;
	assign cst_1_in1_data = forkC_42_out2_data;
	assign cst_1_in1_valid = forkC_42_out2_valid;
	assign forkC_42_out2_ready = cst_1_in1_ready;
	assign cst_2_in1_data = forkC_42_out3_data;
	assign cst_2_in1_valid = forkC_42_out3_valid;
	assign forkC_42_out3_ready = cst_2_in1_ready;
	assign cst_15_in1_data = forkC_42_out4_data;
	assign cst_15_in1_valid = forkC_42_out4_valid;
	assign forkC_42_out4_ready = cst_15_in1_ready;
	assign cst_16_in1_data = forkC_42_out5_data;
	assign cst_16_in1_valid = forkC_42_out5_valid;
	assign forkC_42_out5_ready = cst_16_in1_ready;
	assign branchC_44_in1_data = forkC_42_out6_data;
	assign branchC_44_in1_valid = forkC_42_out6_valid;
	assign forkC_42_out6_ready = branchC_44_in1_ready;
	assign brCst_block1_in1_data = forkC_42_out7_data;
	assign brCst_block1_in1_valid = forkC_42_out7_valid;
	assign forkC_42_out7_ready = brCst_block1_in1_ready;

	assign branchC_44_clk = clk;
	assign branchC_44_rst = rst;
	assign phiC_30_in1_data = branchC_44_out1_data;
	assign phiC_30_in1_valid = branchC_44_out1_valid;
	assign branchC_44_out1_ready = phiC_30_in1_ready;
	assign sink_28_in1_data = branchC_44_out2_data;
	assign sink_28_in1_valid = branchC_44_out2_valid;
	assign branchC_44_out2_ready = sink_28_in1_ready;

	assign brCst_block7_clk = clk;
	assign brCst_block7_rst = rst;
	assign fork_33_in1_data = brCst_block7_out1_data;
	assign fork_33_in1_valid = brCst_block7_out1_valid;
	assign brCst_block7_out1_ready = fork_33_in1_ready;

	assign cst_6_clk = clk;
	assign cst_6_rst = rst;
	assign branch_16_in1_data = cst_6_out1_data;
	assign branch_16_in1_valid = cst_6_out1_valid;
	assign cst_6_out1_ready = branch_16_in1_ready;

	assign cst_7_clk = clk;
	assign cst_7_rst = rst;
	assign branch_17_in1_data = cst_7_out1_data;
	assign branch_17_in1_valid = cst_7_out1_valid;
	assign cst_7_out1_ready = branch_17_in1_ready;

	assign cst_8_clk = clk;
	assign cst_8_rst = rst;
	assign branch_18_in1_data = cst_8_out1_data;
	assign branch_18_in1_valid = cst_8_out1_valid;
	assign cst_8_out1_ready = branch_18_in1_ready;

	assign branch_16_clk = clk;
	assign branch_16_rst = rst;
	assign phi_31_in2_data = branch_16_out1_data;
	assign phi_31_in2_valid = branch_16_out1_valid;
	assign branch_16_out1_ready = phi_31_in2_ready;
	assign sink_12_in1_data = branch_16_out2_data;
	assign sink_12_in1_valid = branch_16_out2_valid;
	assign branch_16_out2_ready = sink_12_in1_ready;

	assign branch_17_clk = clk;
	assign branch_17_rst = rst;
	assign phi_32_in2_data = branch_17_out1_data;
	assign phi_32_in2_valid = branch_17_out1_valid;
	assign branch_17_out1_ready = phi_32_in2_ready;
	assign sink_13_in1_data = branch_17_out2_data;
	assign sink_13_in1_valid = branch_17_out2_valid;
	assign branch_17_out2_ready = sink_13_in1_ready;

	assign branch_18_clk = clk;
	assign branch_18_rst = rst;
	assign phi_33_in2_data = branch_18_out1_data;
	assign phi_33_in2_valid = branch_18_out1_valid;
	assign branch_18_out1_ready = phi_33_in2_ready;
	assign sink_14_in1_data = branch_18_out2_data;
	assign sink_14_in1_valid = branch_18_out2_valid;
	assign branch_18_out2_ready = sink_14_in1_ready;

	assign fork_33_clk = clk;
	assign fork_33_rst = rst;
	assign branch_18_in2_data = fork_33_out1_data;
	assign branch_18_in2_valid = fork_33_out1_valid;
	assign fork_33_out1_ready = branch_18_in2_ready;
	assign branch_17_in2_data = fork_33_out2_data;
	assign branch_17_in2_valid = fork_33_out2_valid;
	assign fork_33_out2_ready = branch_17_in2_ready;
	assign branch_16_in2_data = fork_33_out3_data;
	assign branch_16_in2_valid = fork_33_out3_valid;
	assign fork_33_out3_ready = branch_16_in2_ready;
	assign branchC_50_in2_data = fork_33_out4_data;
	assign branchC_50_in2_valid = fork_33_out4_valid;
	assign fork_33_out4_ready = branchC_50_in2_ready;

	assign phiC_35_clk = clk;
	assign phiC_35_rst = rst;
	assign forkC_48_in1_data = phiC_35_out1_data;
	assign forkC_48_in1_valid = phiC_35_out1_valid;
	assign phiC_35_out1_ready = forkC_48_in1_ready;

	assign forkC_48_clk = clk;
	assign forkC_48_rst = rst;
	assign cst_6_in1_data = forkC_48_out1_data;
	assign cst_6_in1_valid = forkC_48_out1_valid;
	assign forkC_48_out1_ready = cst_6_in1_ready;
	assign cst_7_in1_data = forkC_48_out2_data;
	assign cst_7_in1_valid = forkC_48_out2_valid;
	assign forkC_48_out2_ready = cst_7_in1_ready;
	assign cst_8_in1_data = forkC_48_out3_data;
	assign cst_8_in1_valid = forkC_48_out3_valid;
	assign forkC_48_out3_ready = cst_8_in1_ready;
	assign branchC_50_in1_data = forkC_48_out4_data;
	assign branchC_50_in1_valid = forkC_48_out4_valid;
	assign forkC_48_out4_ready = branchC_50_in1_ready;
	assign brCst_block7_in1_data = forkC_48_out5_data;
	assign brCst_block7_in1_valid = forkC_48_out5_valid;
	assign forkC_48_out5_ready = brCst_block7_in1_ready;

	assign branchC_50_clk = clk;
	assign branchC_50_rst = rst;
	assign phiC_36_in1_data = branchC_50_out1_data;
	assign phiC_36_in1_valid = branchC_50_out1_valid;
	assign branchC_50_out1_ready = phiC_36_in1_ready;
	assign sink_31_in1_data = branchC_50_out2_data;
	assign sink_31_in1_valid = branchC_50_out2_valid;
	assign branchC_50_out2_ready = sink_31_in1_ready;

	assign ret_0_clk = clk;
	assign ret_0_rst = rst;
	assign end_0_in4_data = ret_0_out1_data;
	assign end_0_in4_valid = ret_0_out1_valid;
	assign ret_0_out1_ready = end_0_in4_ready;

	assign phi_n29_clk = clk;
	assign phi_n29_rst = rst;
	assign ret_0_in1_data = phi_n29_out1_data;
	assign ret_0_in1_valid = phi_n29_out1_valid;
	assign phi_n29_out1_ready = ret_0_in1_ready;

	assign end_0_clk = clk;
	assign end_0_rst = rst;
	assign end_out = end_0_out1_data;
	assign end_0_out1_ready = end_ready;
	assign end_valid = end_0_out1_valid;

	assign phiC_43_clk = clk;
	assign phiC_43_rst = rst;
	assign sink_0_in1_data = phiC_43_out1_data;
	assign sink_0_in1_valid = phiC_43_out1_valid;
	assign phiC_43_out1_ready = sink_0_in1_ready;

	assign sink_0_clk = clk;
	assign sink_0_rst = rst;

	assign phi_7_clk = clk;
	assign phi_7_rst = rst;
	assign fork_1_in1_data = phi_7_out1_data;
	assign fork_1_in1_valid = phi_7_out1_valid;
	assign phi_7_out1_ready = fork_1_in1_ready;

	assign cst_3_clk = clk;
	assign cst_3_rst = rst;
	assign icmp_8_in2_data = cst_3_out1_data;
	assign icmp_8_in2_valid = cst_3_out1_valid;
	assign cst_3_out1_ready = icmp_8_in2_ready;

	assign icmp_8_clk = clk;
	assign icmp_8_rst = rst;
	assign fork_29_in1_data = icmp_8_out1_data;
	assign fork_29_in1_valid = icmp_8_out1_valid;
	assign icmp_8_out1_ready = fork_29_in1_ready;

	assign phi_n6_clk = clk;
	assign phi_n6_rst = rst;
	assign branch_6_in1_data = phi_n6_out1_data;
	assign branch_6_in1_valid = phi_n6_out1_valid;
	assign phi_n6_out1_ready = branch_6_in1_ready;

	assign phi_n7_clk = clk;
	assign phi_n7_rst = rst;
	assign branch_7_in1_data = phi_n7_out1_data;
	assign branch_7_in1_valid = phi_n7_out1_valid;
	assign phi_n7_out1_ready = branch_7_in1_ready;

	assign fork_1_clk = clk;
	assign fork_1_rst = rst;
	assign icmp_8_in1_data = fork_1_out1_data;
	assign icmp_8_in1_valid = fork_1_out1_valid;
	assign fork_1_out1_ready = icmp_8_in1_ready;
	assign branch_5_in1_data = fork_1_out2_data;
	assign branch_5_in1_valid = fork_1_out2_valid;
	assign fork_1_out2_ready = branch_5_in1_ready;

	assign branch_5_clk = clk;
	assign branch_5_rst = rst;
	assign phi_n0_in1_data = branch_5_out1_data;
	assign phi_n0_in1_valid = branch_5_out1_valid;
	assign branch_5_out1_ready = phi_n0_in1_ready;
	assign phi_n3_in1_data = branch_5_out2_data;
	assign phi_n3_in1_valid = branch_5_out2_valid;
	assign branch_5_out2_ready = phi_n3_in1_ready;

	assign branch_6_clk = clk;
	assign branch_6_rst = rst;
	assign phi_n1_in1_data = branch_6_out1_data;
	assign phi_n1_in1_valid = branch_6_out1_valid;
	assign branch_6_out1_ready = phi_n1_in1_ready;
	assign phi_n4_in1_data = branch_6_out2_data;
	assign phi_n4_in1_valid = branch_6_out2_valid;
	assign branch_6_out2_ready = phi_n4_in1_ready;

	assign branch_7_clk = clk;
	assign branch_7_rst = rst;
	assign phi_n2_in1_data = branch_7_out1_data;
	assign phi_n2_in1_valid = branch_7_out1_valid;
	assign branch_7_out1_ready = phi_n2_in1_ready;
	assign phi_n5_in1_data = branch_7_out2_data;
	assign phi_n5_in1_valid = branch_7_out2_valid;
	assign branch_7_out2_ready = phi_n5_in1_ready;

	assign fork_29_clk = clk;
	assign fork_29_rst = rst;
	assign branch_7_in2_data = fork_29_out1_data;
	assign branch_7_in2_valid = fork_29_out1_valid;
	assign fork_29_out1_ready = branch_7_in2_ready;
	assign branch_6_in2_data = fork_29_out2_data;
	assign branch_6_in2_valid = fork_29_out2_valid;
	assign fork_29_out2_ready = branch_6_in2_ready;
	assign branch_5_in2_data = fork_29_out3_data;
	assign branch_5_in2_valid = fork_29_out3_valid;
	assign fork_29_out3_ready = branch_5_in2_ready;
	assign branchC_46_in2_data = fork_29_out4_data;
	assign branchC_46_in2_valid = fork_29_out4_valid;
	assign fork_29_out4_ready = branchC_46_in2_ready;

	assign phiC_31_clk = clk;
	assign phiC_31_rst = rst;
	assign branchC_46_in1_data = phiC_31_out1_data;
	assign branchC_46_in1_valid = phiC_31_out1_valid;
	assign phiC_31_out1_ready = branchC_46_in1_ready;
	assign phi_7_in1_data = phiC_31_out2_data;
	assign phi_7_in1_valid = phiC_31_out2_valid;
	assign phiC_31_out2_ready = phi_7_in1_ready;

	assign branchC_46_clk = clk;
	assign branchC_46_rst = rst;
	assign phiC_32_in1_data = branchC_46_out1_data;
	assign phiC_32_in1_valid = branchC_46_out1_valid;
	assign branchC_46_out1_ready = phiC_32_in1_ready;
	assign phiC_34_in1_data = branchC_46_out2_data;
	assign phiC_34_in1_valid = branchC_46_out2_valid;
	assign branchC_46_out2_ready = phiC_34_in1_ready;

	assign source_0_clk = clk;
	assign source_0_rst = rst;
	assign cst_3_in1_data = source_0_out1_data;
	assign cst_3_in1_valid = source_0_out1_valid;
	assign source_0_out1_ready = cst_3_in1_ready;

	assign load_17_clk = clk;
	assign load_17_rst = rst;
	assign branch_11_in1_data = load_17_out1_data;
	assign branch_11_in1_valid = load_17_out1_valid;
	assign load_17_out1_ready = branch_11_in1_ready;
	assign MC_kmpNext_in5_data = load_17_out2_data;
	assign MC_kmpNext_in5_valid = load_17_out2_valid;
	assign load_17_out2_ready = MC_kmpNext_in5_ready;

	assign brCst_block5_clk = clk;
	assign brCst_block5_rst = rst;
	assign fork_31_in1_data = brCst_block5_out1_data;
	assign fork_31_in1_valid = brCst_block5_out1_valid;
	assign brCst_block5_out1_ready = fork_31_in1_ready;

	assign phi_n8_clk = clk;
	assign phi_n8_rst = rst;
	assign fork_16_in1_data = phi_n8_out1_data;
	assign fork_16_in1_valid = phi_n8_out1_valid;
	assign phi_n8_out1_ready = fork_16_in1_ready;

	assign phi_n9_clk = clk;
	assign phi_n9_rst = rst;
	assign branch_12_in1_data = phi_n9_out1_data;
	assign branch_12_in1_valid = phi_n9_out1_valid;
	assign phi_n9_out1_ready = branch_12_in1_ready;

	assign fork_16_clk = clk;
	assign fork_16_rst = rst;
	assign load_17_in2_data = fork_16_out1_data;
	assign load_17_in2_valid = fork_16_out1_valid;
	assign fork_16_out1_ready = load_17_in2_ready;
	assign branch_13_in1_data = fork_16_out2_data;
	assign branch_13_in1_valid = fork_16_out2_valid;
	assign fork_16_out2_ready = branch_13_in1_ready;

	assign branch_11_clk = clk;
	assign branch_11_rst = rst;
	assign Buffer_100_in1_data = branch_11_out1_data;
	assign Buffer_100_in1_valid = branch_11_out1_valid;
	assign branch_11_out1_ready = Buffer_100_in1_ready;
	assign sink_7_in1_data = branch_11_out2_data;
	assign sink_7_in1_valid = branch_11_out2_valid;
	assign branch_11_out2_ready = sink_7_in1_ready;

	assign branch_12_clk = clk;
	assign branch_12_rst = rst;
	assign Buffer_101_in1_data = branch_12_out1_data;
	assign Buffer_101_in1_valid = branch_12_out1_valid;
	assign branch_12_out1_ready = Buffer_101_in1_ready;
	assign sink_8_in1_data = branch_12_out2_data;
	assign sink_8_in1_valid = branch_12_out2_valid;
	assign branch_12_out2_ready = sink_8_in1_ready;

	assign branch_13_clk = clk;
	assign branch_13_rst = rst;
	assign Buffer_102_in1_data = branch_13_out1_data;
	assign Buffer_102_in1_valid = branch_13_out1_valid;
	assign branch_13_out1_ready = Buffer_102_in1_ready;
	assign sink_9_in1_data = branch_13_out2_data;
	assign sink_9_in1_valid = branch_13_out2_valid;
	assign branch_13_out2_ready = sink_9_in1_ready;

	assign fork_31_clk = clk;
	assign fork_31_rst = rst;
	assign branch_13_in2_data = fork_31_out1_data;
	assign branch_13_in2_valid = fork_31_out1_valid;
	assign fork_31_out1_ready = branch_13_in2_ready;
	assign branch_12_in2_data = fork_31_out2_data;
	assign branch_12_in2_valid = fork_31_out2_valid;
	assign fork_31_out2_ready = branch_12_in2_ready;
	assign branch_11_in2_data = fork_31_out3_data;
	assign branch_11_in2_valid = fork_31_out3_valid;
	assign fork_31_out3_ready = branch_11_in2_ready;
	assign branchC_48_in2_data = fork_31_out4_data;
	assign branchC_48_in2_valid = fork_31_out4_valid;
	assign fork_31_out4_ready = branchC_48_in2_ready;

	assign phiC_33_clk = clk;
	assign phiC_33_rst = rst;
	assign forkC_46_in1_data = phiC_33_out1_data;
	assign forkC_46_in1_valid = phiC_33_out1_valid;
	assign phiC_33_out1_ready = forkC_46_in1_ready;

	assign forkC_46_clk = clk;
	assign forkC_46_rst = rst;
	assign branchC_48_in1_data = forkC_46_out1_data;
	assign branchC_48_in1_valid = forkC_46_out1_valid;
	assign forkC_46_out1_ready = branchC_48_in1_ready;
	assign brCst_block5_in1_data = forkC_46_out2_data;
	assign brCst_block5_in1_valid = forkC_46_out2_valid;
	assign forkC_46_out2_ready = brCst_block5_in1_ready;

	assign branchC_48_clk = clk;
	assign branchC_48_rst = rst;
	assign Buffer_103_in1_data = branchC_48_out1_data;
	assign Buffer_103_in1_valid = branchC_48_out1_valid;
	assign branchC_48_out1_ready = Buffer_103_in1_ready;
	assign sink_30_in1_data = branchC_48_out2_data;
	assign sink_30_in1_valid = branchC_48_out2_valid;
	assign branchC_48_out2_ready = sink_30_in1_ready;

	assign phi_38_clk = clk;
	assign phi_38_rst = rst;
	assign fork_5_in1_data = phi_38_out1_data;
	assign fork_5_in1_valid = phi_38_out1_valid;
	assign phi_38_out1_ready = fork_5_in1_ready;

	assign cst_9_clk = clk;
	assign cst_9_rst = rst;
	assign icmp_39_in2_data = cst_9_out1_data;
	assign icmp_39_in2_valid = cst_9_out1_valid;
	assign cst_9_out1_ready = icmp_39_in2_ready;

	assign icmp_39_clk = clk;
	assign icmp_39_rst = rst;
	assign fork_35_in1_data = icmp_39_out1_data;
	assign fork_35_in1_valid = icmp_39_out1_valid;
	assign icmp_39_out1_ready = fork_35_in1_ready;

	assign phi_n10_clk = clk;
	assign phi_n10_rst = rst;
	assign branch_24_in1_data = phi_n10_out1_data;
	assign branch_24_in1_valid = phi_n10_out1_valid;
	assign phi_n10_out1_ready = branch_24_in1_ready;

	assign phi_n11_clk = clk;
	assign phi_n11_rst = rst;
	assign branch_25_in1_data = phi_n11_out1_data;
	assign branch_25_in1_valid = phi_n11_out1_valid;
	assign phi_n11_out1_ready = branch_25_in1_ready;

	assign phi_n12_clk = clk;
	assign phi_n12_rst = rst;
	assign branch_26_in1_data = phi_n12_out1_data;
	assign branch_26_in1_valid = phi_n12_out1_valid;
	assign phi_n12_out1_ready = branch_26_in1_ready;

	assign fork_5_clk = clk;
	assign fork_5_rst = rst;
	assign icmp_39_in1_data = fork_5_out1_data;
	assign icmp_39_in1_valid = fork_5_out1_valid;
	assign fork_5_out1_ready = icmp_39_in1_ready;
	assign branch_23_in1_data = fork_5_out2_data;
	assign branch_23_in1_valid = fork_5_out2_valid;
	assign fork_5_out2_ready = branch_23_in1_ready;

	assign branch_23_clk = clk;
	assign branch_23_rst = rst;
	assign phi_n21_in1_data = branch_23_out1_data;
	assign phi_n21_in1_valid = branch_23_out1_valid;
	assign branch_23_out1_ready = phi_n21_in1_ready;
	assign phi_n25_in1_data = branch_23_out2_data;
	assign phi_n25_in1_valid = branch_23_out2_valid;
	assign branch_23_out2_ready = phi_n25_in1_ready;

	assign branch_24_clk = clk;
	assign branch_24_rst = rst;
	assign phi_n22_in1_data = branch_24_out1_data;
	assign phi_n22_in1_valid = branch_24_out1_valid;
	assign branch_24_out1_ready = phi_n22_in1_ready;
	assign phi_n26_in1_data = branch_24_out2_data;
	assign phi_n26_in1_valid = branch_24_out2_valid;
	assign branch_24_out2_ready = phi_n26_in1_ready;

	assign branch_25_clk = clk;
	assign branch_25_rst = rst;
	assign phi_n23_in1_data = branch_25_out1_data;
	assign phi_n23_in1_valid = branch_25_out1_valid;
	assign branch_25_out1_ready = phi_n23_in1_ready;
	assign phi_n27_in1_data = branch_25_out2_data;
	assign phi_n27_in1_valid = branch_25_out2_valid;
	assign branch_25_out2_ready = phi_n27_in1_ready;

	assign branch_26_clk = clk;
	assign branch_26_rst = rst;
	assign phi_n24_in1_data = branch_26_out1_data;
	assign phi_n24_in1_valid = branch_26_out1_valid;
	assign branch_26_out1_ready = phi_n24_in1_ready;
	assign phi_n28_in1_data = branch_26_out2_data;
	assign phi_n28_in1_valid = branch_26_out2_valid;
	assign branch_26_out2_ready = phi_n28_in1_ready;

	assign fork_35_clk = clk;
	assign fork_35_rst = rst;
	assign branch_26_in2_data = fork_35_out1_data;
	assign branch_26_in2_valid = fork_35_out1_valid;
	assign fork_35_out1_ready = branch_26_in2_ready;
	assign branch_25_in2_data = fork_35_out2_data;
	assign branch_25_in2_valid = fork_35_out2_valid;
	assign fork_35_out2_ready = branch_25_in2_ready;
	assign branch_24_in2_data = fork_35_out3_data;
	assign branch_24_in2_valid = fork_35_out3_valid;
	assign fork_35_out3_ready = branch_24_in2_ready;
	assign branch_23_in2_data = fork_35_out4_data;
	assign branch_23_in2_valid = fork_35_out4_valid;
	assign fork_35_out4_ready = branch_23_in2_ready;
	assign branchC_52_in2_data = fork_35_out5_data;
	assign branchC_52_in2_valid = fork_35_out5_valid;
	assign fork_35_out5_ready = branchC_52_in2_ready;

	assign phiC_37_clk = clk;
	assign phiC_37_rst = rst;
	assign branchC_52_in1_data = phiC_37_out1_data;
	assign branchC_52_in1_valid = phiC_37_out1_valid;
	assign phiC_37_out1_ready = branchC_52_in1_ready;
	assign phi_38_in1_data = phiC_37_out2_data;
	assign phi_38_in1_valid = phiC_37_out2_valid;
	assign phiC_37_out2_ready = phi_38_in1_ready;

	assign branchC_52_clk = clk;
	assign branchC_52_rst = rst;
	assign phiC_38_in1_data = branchC_52_out1_data;
	assign phiC_38_in1_valid = branchC_52_out1_valid;
	assign branchC_52_out1_ready = phiC_38_in1_ready;
	assign phiC_40_in1_data = branchC_52_out2_data;
	assign phiC_40_in1_valid = branchC_52_out2_valid;
	assign branchC_52_out2_ready = phiC_40_in1_ready;

	assign source_3_clk = clk;
	assign source_3_rst = rst;
	assign cst_9_in1_data = source_3_out1_data;
	assign cst_9_in1_valid = source_3_out1_valid;
	assign source_3_out1_ready = cst_9_in1_ready;

	assign load_21_clk = clk;
	assign load_21_rst = rst;
	assign icmp_22_in1_data = load_21_out1_data;
	assign icmp_22_in1_valid = load_21_out1_valid;
	assign load_21_out1_ready = icmp_22_in1_ready;
	assign MC_pattern_in3_data = load_21_out2_data;
	assign MC_pattern_in3_valid = load_21_out2_valid;
	assign load_21_out2_ready = MC_pattern_in3_ready;

	assign icmp_22_clk = clk;
	assign icmp_22_rst = rst;
	assign zext_23_in1_data = icmp_22_out1_data;
	assign zext_23_in1_valid = icmp_22_out1_valid;
	assign icmp_22_out1_ready = zext_23_in1_ready;

	assign zext_23_clk = clk;
	assign zext_23_rst = rst;
	assign add_24_in2_data = zext_23_out1_data;
	assign add_24_in2_valid = zext_23_out1_valid;
	assign zext_23_out1_ready = add_24_in2_ready;

	assign add_24_clk = clk;
	assign add_24_rst = rst;
	assign fork_2_in1_data = add_24_out1_data;
	assign fork_2_in1_valid = add_24_out1_valid;
	assign add_24_out1_ready = fork_2_in1_ready;

	assign store_1_clk = clk;
	assign store_1_rst = rst;
	assign MC_kmpNext_in7_data = store_1_out1_data;
	assign MC_kmpNext_in7_valid = store_1_out1_valid;
	assign store_1_out1_ready = MC_kmpNext_in7_ready;
	assign MC_kmpNext_in6_data = store_1_out2_data;
	assign MC_kmpNext_in6_valid = store_1_out2_valid;
	assign store_1_out2_ready = MC_kmpNext_in6_ready;

	assign cst_4_clk = clk;
	assign cst_4_rst = rst;
	assign add_27_in2_data = cst_4_out1_data;
	assign add_27_in2_valid = cst_4_out1_valid;
	assign cst_4_out1_ready = add_27_in2_ready;

	assign add_27_clk = clk;
	assign add_27_rst = rst;
	assign fork_3_in1_data = add_27_out1_data;
	assign fork_3_in1_valid = add_27_out1_valid;
	assign add_27_out1_ready = fork_3_in1_ready;

	assign cst_5_clk = clk;
	assign cst_5_rst = rst;
	assign icmp_28_in2_data = cst_5_out1_data;
	assign icmp_28_in2_valid = cst_5_out1_valid;
	assign cst_5_out1_ready = icmp_28_in2_ready;

	assign icmp_28_clk = clk;
	assign icmp_28_rst = rst;
	assign fork_32_in1_data = icmp_28_out1_data;
	assign fork_32_in1_valid = icmp_28_out1_valid;
	assign icmp_28_out1_ready = fork_32_in1_ready;

	assign phi_n3_clk = clk;
	assign phi_n3_rst = rst;
	assign fork_12_in1_data = phi_n3_out1_data;
	assign fork_12_in1_valid = phi_n3_out1_valid;
	assign phi_n3_out1_ready = fork_12_in1_ready;

	assign phi_n4_clk = clk;
	assign phi_n4_rst = rst;
	assign icmp_22_in2_data = phi_n4_out1_data;
	assign icmp_22_in2_valid = phi_n4_out1_valid;
	assign phi_n4_out1_ready = icmp_22_in2_ready;

	assign phi_n5_clk = clk;
	assign phi_n5_rst = rst;
	assign fork_13_in1_data = phi_n5_out1_data;
	assign fork_13_in1_valid = phi_n5_out1_valid;
	assign phi_n5_out1_ready = fork_13_in1_ready;

	assign fork_2_clk = clk;
	assign fork_2_rst = rst;
	assign store_1_in1_data = fork_2_out1_data;
	assign store_1_in1_valid = fork_2_out1_valid;
	assign fork_2_out1_ready = store_1_in1_ready;
	assign branch_14_in1_data = fork_2_out2_data;
	assign branch_14_in1_valid = fork_2_out2_valid;
	assign fork_2_out2_ready = branch_14_in1_ready;

	assign fork_3_clk = clk;
	assign fork_3_rst = rst;
	assign icmp_28_in1_data = fork_3_out1_data;
	assign icmp_28_in1_valid = fork_3_out1_valid;
	assign fork_3_out1_ready = icmp_28_in1_ready;
	assign branch_15_in1_data = fork_3_out2_data;
	assign branch_15_in1_valid = fork_3_out2_valid;
	assign fork_3_out2_ready = branch_15_in1_ready;

	assign fork_12_clk = clk;
	assign fork_12_rst = rst;
	assign load_21_in2_data = fork_12_out1_data;
	assign load_21_in2_valid = fork_12_out1_valid;
	assign fork_12_out1_ready = load_21_in2_ready;
	assign add_24_in1_data = fork_12_out2_data;
	assign add_24_in1_valid = fork_12_out2_valid;
	assign fork_12_out2_ready = add_24_in1_ready;

	assign fork_13_clk = clk;
	assign fork_13_rst = rst;
	assign store_1_in2_data = fork_13_out1_data;
	assign store_1_in2_valid = fork_13_out1_valid;
	assign fork_13_out1_ready = store_1_in2_ready;
	assign add_27_in1_data = fork_13_out2_data;
	assign add_27_in1_valid = fork_13_out2_valid;
	assign fork_13_out2_ready = add_27_in1_ready;

	assign branch_14_clk = clk;
	assign branch_14_rst = rst;
	assign Buffer_104_in1_data = branch_14_out1_data;
	assign Buffer_104_in1_valid = branch_14_out1_valid;
	assign branch_14_out1_ready = Buffer_104_in1_ready;
	assign sink_10_in1_data = branch_14_out2_data;
	assign sink_10_in1_valid = branch_14_out2_valid;
	assign branch_14_out2_ready = sink_10_in1_ready;

	assign branch_15_clk = clk;
	assign branch_15_rst = rst;
	assign Buffer_105_in1_data = branch_15_out1_data;
	assign Buffer_105_in1_valid = branch_15_out1_valid;
	assign branch_15_out1_ready = Buffer_105_in1_ready;
	assign sink_11_in1_data = branch_15_out2_data;
	assign sink_11_in1_valid = branch_15_out2_valid;
	assign branch_15_out2_ready = sink_11_in1_ready;

	assign fork_32_clk = clk;
	assign fork_32_rst = rst;
	assign branch_15_in2_data = fork_32_out1_data;
	assign branch_15_in2_valid = fork_32_out1_valid;
	assign fork_32_out1_ready = branch_15_in2_ready;
	assign branch_14_in2_data = fork_32_out2_data;
	assign branch_14_in2_valid = fork_32_out2_valid;
	assign fork_32_out2_ready = branch_14_in2_ready;
	assign branchC_49_in2_data = fork_32_out3_data;
	assign branchC_49_in2_valid = fork_32_out3_valid;
	assign fork_32_out3_ready = branchC_49_in2_ready;

	assign cst_17_clk = clk;
	assign cst_17_rst = rst;
	assign MC_kmpNext_in2_data = cst_17_out1_data;
	assign MC_kmpNext_in2_valid = cst_17_out1_valid;
	assign cst_17_out1_ready = MC_kmpNext_in2_ready;

	assign phiC_34_clk = clk;
	assign phiC_34_rst = rst;
	assign forkC_47_in1_data = phiC_34_out1_data;
	assign forkC_47_in1_valid = phiC_34_out1_valid;
	assign phiC_34_out1_ready = forkC_47_in1_ready;

	assign forkC_47_clk = clk;
	assign forkC_47_rst = rst;
	assign cst_17_in1_data = forkC_47_out1_data;
	assign cst_17_in1_valid = forkC_47_out1_valid;
	assign forkC_47_out1_ready = cst_17_in1_ready;
	assign branchC_49_in1_data = forkC_47_out2_data;
	assign branchC_49_in1_valid = forkC_47_out2_valid;
	assign forkC_47_out2_ready = branchC_49_in1_ready;

	assign branchC_49_clk = clk;
	assign branchC_49_rst = rst;
	assign Buffer_106_in1_data = branchC_49_out1_data;
	assign Buffer_106_in1_valid = branchC_49_out1_valid;
	assign branchC_49_out1_ready = Buffer_106_in1_ready;
	assign phiC_35_in1_data = branchC_49_out2_data;
	assign phiC_35_in1_valid = branchC_49_out2_valid;
	assign branchC_49_out2_ready = phiC_35_in1_ready;

	assign source_1_clk = clk;
	assign source_1_rst = rst;
	assign cst_4_in1_data = source_1_out1_data;
	assign cst_4_in1_valid = source_1_out1_valid;
	assign source_1_out1_ready = cst_4_in1_ready;

	assign source_2_clk = clk;
	assign source_2_rst = rst;
	assign cst_5_in1_data = source_2_out1_data;
	assign cst_5_in1_valid = source_2_out1_valid;
	assign source_2_out1_ready = cst_5_in1_ready;

	assign load_12_clk = clk;
	assign load_12_rst = rst;
	assign icmp_13_in1_data = load_12_out1_data;
	assign icmp_13_in1_valid = load_12_out1_valid;
	assign load_12_out1_ready = icmp_13_in1_ready;
	assign MC_pattern_in2_data = load_12_out2_data;
	assign MC_pattern_in2_valid = load_12_out2_valid;
	assign load_12_out2_ready = MC_pattern_in2_ready;

	assign icmp_13_clk = clk;
	assign icmp_13_rst = rst;
	assign fork_30_in1_data = icmp_13_out1_data;
	assign fork_30_in1_valid = icmp_13_out1_valid;
	assign icmp_13_out1_ready = fork_30_in1_ready;

	assign phi_n0_clk = clk;
	assign phi_n0_rst = rst;
	assign fork_9_in1_data = phi_n0_out1_data;
	assign fork_9_in1_valid = phi_n0_out1_valid;
	assign phi_n0_out1_ready = fork_9_in1_ready;

	assign phi_n1_clk = clk;
	assign phi_n1_rst = rst;
	assign fork_10_in1_data = phi_n1_out1_data;
	assign fork_10_in1_valid = phi_n1_out1_valid;
	assign phi_n1_out1_ready = fork_10_in1_ready;

	assign phi_n2_clk = clk;
	assign phi_n2_rst = rst;
	assign branch_10_in1_data = phi_n2_out1_data;
	assign branch_10_in1_valid = phi_n2_out1_valid;
	assign phi_n2_out1_ready = branch_10_in1_ready;

	assign fork_9_clk = clk;
	assign fork_9_rst = rst;
	assign load_12_in2_data = fork_9_out1_data;
	assign load_12_in2_valid = fork_9_out1_valid;
	assign fork_9_out1_ready = load_12_in2_ready;
	assign branch_8_in1_data = fork_9_out2_data;
	assign branch_8_in1_valid = fork_9_out2_valid;
	assign fork_9_out2_ready = branch_8_in1_ready;

	assign fork_10_clk = clk;
	assign fork_10_rst = rst;
	assign icmp_13_in2_data = fork_10_out1_data;
	assign icmp_13_in2_valid = fork_10_out1_valid;
	assign fork_10_out1_ready = icmp_13_in2_ready;
	assign branch_9_in1_data = fork_10_out2_data;
	assign branch_9_in1_valid = fork_10_out2_valid;
	assign fork_10_out2_ready = branch_9_in1_ready;

	assign branch_8_clk = clk;
	assign branch_8_rst = rst;
	assign phi_n3_in2_data = branch_8_out1_data;
	assign phi_n3_in2_valid = branch_8_out1_valid;
	assign branch_8_out1_ready = phi_n3_in2_ready;
	assign sink_6_in1_data = branch_8_out2_data;
	assign sink_6_in1_valid = branch_8_out2_valid;
	assign branch_8_out2_ready = sink_6_in1_ready;

	assign branch_9_clk = clk;
	assign branch_9_rst = rst;
	assign phi_n4_in2_data = branch_9_out1_data;
	assign phi_n4_in2_valid = branch_9_out1_valid;
	assign branch_9_out1_ready = phi_n4_in2_ready;
	assign phi_n9_in1_data = branch_9_out2_data;
	assign phi_n9_in1_valid = branch_9_out2_valid;
	assign branch_9_out2_ready = phi_n9_in1_ready;

	assign branch_10_clk = clk;
	assign branch_10_rst = rst;
	assign phi_n5_in2_data = branch_10_out1_data;
	assign phi_n5_in2_valid = branch_10_out1_valid;
	assign branch_10_out1_ready = phi_n5_in2_ready;
	assign phi_n8_in1_data = branch_10_out2_data;
	assign phi_n8_in1_valid = branch_10_out2_valid;
	assign branch_10_out2_ready = phi_n8_in1_ready;

	assign fork_30_clk = clk;
	assign fork_30_rst = rst;
	assign branch_10_in2_data = fork_30_out1_data;
	assign branch_10_in2_valid = fork_30_out1_valid;
	assign fork_30_out1_ready = branch_10_in2_ready;
	assign branch_9_in2_data = fork_30_out2_data;
	assign branch_9_in2_valid = fork_30_out2_valid;
	assign fork_30_out2_ready = branch_9_in2_ready;
	assign branch_8_in2_data = fork_30_out3_data;
	assign branch_8_in2_valid = fork_30_out3_valid;
	assign fork_30_out3_ready = branch_8_in2_ready;
	assign branchC_47_in2_data = fork_30_out4_data;
	assign branchC_47_in2_valid = fork_30_out4_valid;
	assign fork_30_out4_ready = branchC_47_in2_ready;

	assign phiC_32_clk = clk;
	assign phiC_32_rst = rst;
	assign branchC_47_in1_data = phiC_32_out1_data;
	assign branchC_47_in1_valid = phiC_32_out1_valid;
	assign phiC_32_out1_ready = branchC_47_in1_ready;

	assign branchC_47_clk = clk;
	assign branchC_47_rst = rst;
	assign phiC_34_in2_data = branchC_47_out1_data;
	assign phiC_34_in2_valid = branchC_47_out1_valid;
	assign branchC_47_out1_ready = phiC_34_in2_ready;
	assign phiC_33_in1_data = branchC_47_out2_data;
	assign phiC_33_in1_valid = branchC_47_out2_valid;
	assign branchC_47_out2_ready = phiC_33_in1_ready;

	assign phi_64_clk = clk;
	assign phi_64_rst = rst;
	assign branch_41_in1_data = phi_64_out1_data;
	assign branch_41_in1_valid = phi_64_out1_valid;
	assign phi_64_out1_ready = branch_41_in1_ready;

	assign phi_65_clk = clk;
	assign phi_65_rst = rst;
	assign branch_42_in1_data = phi_65_out1_data;
	assign branch_42_in1_valid = phi_65_out1_valid;
	assign phi_65_out1_ready = branch_42_in1_ready;

	assign cst_13_clk = clk;
	assign cst_13_rst = rst;
	assign add_66_in2_data = cst_13_out1_data;
	assign add_66_in2_valid = cst_13_out1_valid;
	assign cst_13_out1_ready = add_66_in2_ready;

	assign add_66_clk = clk;
	assign add_66_rst = rst;
	assign fork_8_in1_data = add_66_out1_data;
	assign fork_8_in1_valid = add_66_out1_valid;
	assign add_66_out1_ready = fork_8_in1_ready;

	assign cst_14_clk = clk;
	assign cst_14_rst = rst;
	assign icmp_67_in2_data = cst_14_out1_data;
	assign icmp_67_in2_valid = cst_14_out1_valid;
	assign cst_14_out1_ready = icmp_67_in2_ready;

	assign icmp_67_clk = clk;
	assign icmp_67_rst = rst;
	assign fork_40_in1_data = icmp_67_out1_data;
	assign fork_40_in1_valid = icmp_67_out1_valid;
	assign icmp_67_out1_ready = fork_40_in1_ready;

	assign phi_n16_clk = clk;
	assign phi_n16_rst = rst;
	assign add_66_in1_data = phi_n16_out1_data;
	assign add_66_in1_valid = phi_n16_out1_valid;
	assign phi_n16_out1_ready = add_66_in1_ready;

	assign fork_8_clk = clk;
	assign fork_8_rst = rst;
	assign icmp_67_in1_data = fork_8_out1_data;
	assign icmp_67_in1_valid = fork_8_out1_valid;
	assign fork_8_out1_ready = icmp_67_in1_ready;
	assign branch_43_in1_data = fork_8_out2_data;
	assign branch_43_in1_valid = fork_8_out2_valid;
	assign fork_8_out2_ready = branch_43_in1_ready;

	assign branch_41_clk = clk;
	assign branch_41_rst = rst;
	assign Buffer_112_in1_data = branch_41_out1_data;
	assign Buffer_112_in1_valid = branch_41_out1_valid;
	assign branch_41_out1_ready = Buffer_112_in1_ready;
	assign sink_26_in1_data = branch_41_out2_data;
	assign sink_26_in1_valid = branch_41_out2_valid;
	assign branch_41_out2_ready = sink_26_in1_ready;

	assign branch_42_clk = clk;
	assign branch_42_rst = rst;
	assign Buffer_113_in1_data = branch_42_out1_data;
	assign Buffer_113_in1_valid = branch_42_out1_valid;
	assign branch_42_out1_ready = Buffer_113_in1_ready;
	assign phi_n29_in1_data = branch_42_out2_data;
	assign phi_n29_in1_valid = branch_42_out2_valid;
	assign branch_42_out2_ready = phi_n29_in1_ready;

	assign branch_43_clk = clk;
	assign branch_43_rst = rst;
	assign Buffer_114_in1_data = branch_43_out1_data;
	assign Buffer_114_in1_valid = branch_43_out1_valid;
	assign branch_43_out1_ready = Buffer_114_in1_ready;
	assign sink_27_in1_data = branch_43_out2_data;
	assign sink_27_in1_valid = branch_43_out2_valid;
	assign branch_43_out2_ready = sink_27_in1_ready;

	assign fork_40_clk = clk;
	assign fork_40_rst = rst;
	assign branch_43_in2_data = fork_40_out1_data;
	assign branch_43_in2_valid = fork_40_out1_valid;
	assign fork_40_out1_ready = branch_43_in2_ready;
	assign branch_42_in2_data = fork_40_out2_data;
	assign branch_42_in2_valid = fork_40_out2_valid;
	assign fork_40_out2_ready = branch_42_in2_ready;
	assign branch_41_in2_data = fork_40_out3_data;
	assign branch_41_in2_valid = fork_40_out3_valid;
	assign fork_40_out3_ready = branch_41_in2_ready;
	assign branchC_57_in2_data = fork_40_out4_data;
	assign branchC_57_in2_valid = fork_40_out4_valid;
	assign fork_40_out4_ready = branchC_57_in2_ready;

	assign phiC_42_clk = clk;
	assign phiC_42_rst = rst;
	assign branchC_57_in1_data = phiC_42_out1_data;
	assign branchC_57_in1_valid = phiC_42_out1_valid;
	assign phiC_42_out1_ready = branchC_57_in1_ready;
	assign fork_61_in1_data = phiC_42_out2_data;
	assign fork_61_in1_valid = phiC_42_out2_valid;
	assign phiC_42_out2_ready = fork_61_in1_ready;

	assign branchC_57_clk = clk;
	assign branchC_57_rst = rst;
	assign Buffer_115_in1_data = branchC_57_out1_data;
	assign Buffer_115_in1_valid = branchC_57_out1_valid;
	assign branchC_57_out1_ready = Buffer_115_in1_ready;
	assign phiC_43_in1_data = branchC_57_out2_data;
	assign phiC_43_in1_valid = branchC_57_out2_valid;
	assign branchC_57_out2_ready = phiC_43_in1_ready;

	assign source_7_clk = clk;
	assign source_7_rst = rst;
	assign cst_13_in1_data = source_7_out1_data;
	assign cst_13_in1_valid = source_7_out1_valid;
	assign source_7_out1_ready = cst_13_in1_ready;

	assign source_8_clk = clk;
	assign source_8_rst = rst;
	assign cst_14_in1_data = source_8_out1_data;
	assign cst_14_in1_valid = source_8_out1_valid;
	assign source_8_out1_ready = cst_14_in1_ready;

	assign fork_61_clk = clk;
	assign fork_61_rst = rst;
	assign phi_64_in1_data = fork_61_out1_data;
	assign phi_64_in1_valid = fork_61_out1_valid;
	assign fork_61_out1_ready = phi_64_in1_ready;
	assign phi_65_in1_data = fork_61_out2_data;
	assign phi_65_in1_valid = fork_61_out2_valid;
	assign fork_61_out2_ready = phi_65_in1_ready;

	assign cst_11_clk = clk;
	assign cst_11_rst = rst;
	assign add_58_in2_data = cst_11_out1_data;
	assign add_58_in2_valid = cst_11_out1_valid;
	assign cst_11_out1_ready = add_58_in2_ready;

	assign add_58_clk = clk;
	assign add_58_rst = rst;
	assign branch_39_in1_data = add_58_out1_data;
	assign branch_39_in1_valid = add_58_out1_valid;
	assign add_58_out1_ready = branch_39_in1_ready;

	assign cst_12_clk = clk;
	assign cst_12_rst = rst;
	assign add_59_in2_data = cst_12_out1_data;
	assign add_59_in2_valid = cst_12_out1_valid;
	assign cst_12_out1_ready = add_59_in2_ready;

	assign add_59_clk = clk;
	assign add_59_rst = rst;
	assign load_62_in2_data = add_59_out1_data;
	assign load_62_in2_valid = add_59_out1_valid;
	assign add_59_out1_ready = load_62_in2_ready;

	assign load_62_clk = clk;
	assign load_62_rst = rst;
	assign branch_38_in1_data = load_62_out1_data;
	assign branch_38_in1_valid = load_62_out1_valid;
	assign load_62_out1_ready = branch_38_in1_ready;
	assign MC_kmpNext_in9_data = load_62_out2_data;
	assign MC_kmpNext_in9_valid = load_62_out2_valid;
	assign load_62_out2_ready = MC_kmpNext_in9_ready;

	assign brCst_block13_clk = clk;
	assign brCst_block13_rst = rst;
	assign fork_39_in1_data = brCst_block13_out1_data;
	assign fork_39_in1_valid = brCst_block13_out1_valid;
	assign brCst_block13_out1_ready = fork_39_in1_ready;

	assign phi_n13_clk = clk;
	assign phi_n13_rst = rst;
	assign add_58_in1_data = phi_n13_out1_data;
	assign add_58_in1_valid = phi_n13_out1_valid;
	assign phi_n13_out1_ready = add_58_in1_ready;

	assign phi_n14_clk = clk;
	assign phi_n14_rst = rst;
	assign add_59_in1_data = phi_n14_out1_data;
	assign add_59_in1_valid = phi_n14_out1_valid;
	assign phi_n14_out1_ready = add_59_in1_ready;

	assign phi_n15_clk = clk;
	assign phi_n15_rst = rst;
	assign branch_40_in1_data = phi_n15_out1_data;
	assign branch_40_in1_valid = phi_n15_out1_valid;
	assign phi_n15_out1_ready = branch_40_in1_ready;

	assign branch_38_clk = clk;
	assign branch_38_rst = rst;
	assign phi_64_in3_data = branch_38_out1_data;
	assign phi_64_in3_valid = branch_38_out1_valid;
	assign branch_38_out1_ready = phi_64_in3_ready;
	assign sink_23_in1_data = branch_38_out2_data;
	assign sink_23_in1_valid = branch_38_out2_valid;
	assign branch_38_out2_ready = sink_23_in1_ready;

	assign branch_39_clk = clk;
	assign branch_39_rst = rst;
	assign phi_65_in3_data = branch_39_out1_data;
	assign phi_65_in3_valid = branch_39_out1_valid;
	assign branch_39_out1_ready = phi_65_in3_ready;
	assign sink_24_in1_data = branch_39_out2_data;
	assign sink_24_in1_valid = branch_39_out2_valid;
	assign branch_39_out2_ready = sink_24_in1_ready;

	assign branch_40_clk = clk;
	assign branch_40_rst = rst;
	assign phi_n16_in2_data = branch_40_out1_data;
	assign phi_n16_in2_valid = branch_40_out1_valid;
	assign branch_40_out1_ready = phi_n16_in2_ready;
	assign sink_25_in1_data = branch_40_out2_data;
	assign sink_25_in1_valid = branch_40_out2_valid;
	assign branch_40_out2_ready = sink_25_in1_ready;

	assign fork_39_clk = clk;
	assign fork_39_rst = rst;
	assign branch_40_in2_data = fork_39_out1_data;
	assign branch_40_in2_valid = fork_39_out1_valid;
	assign fork_39_out1_ready = branch_40_in2_ready;
	assign branch_39_in2_data = fork_39_out2_data;
	assign branch_39_in2_valid = fork_39_out2_valid;
	assign fork_39_out2_ready = branch_39_in2_ready;
	assign branch_38_in2_data = fork_39_out3_data;
	assign branch_38_in2_valid = fork_39_out3_valid;
	assign fork_39_out3_ready = branch_38_in2_ready;
	assign branchC_56_in2_data = fork_39_out4_data;
	assign branchC_56_in2_valid = fork_39_out4_valid;
	assign fork_39_out4_ready = branchC_56_in2_ready;

	assign phiC_41_clk = clk;
	assign phiC_41_rst = rst;
	assign forkC_54_in1_data = phiC_41_out1_data;
	assign forkC_54_in1_valid = phiC_41_out1_valid;
	assign phiC_41_out1_ready = forkC_54_in1_ready;

	assign forkC_54_clk = clk;
	assign forkC_54_rst = rst;
	assign branchC_56_in1_data = forkC_54_out1_data;
	assign branchC_56_in1_valid = forkC_54_out1_valid;
	assign forkC_54_out1_ready = branchC_56_in1_ready;
	assign brCst_block13_in1_data = forkC_54_out2_data;
	assign brCst_block13_in1_valid = forkC_54_out2_valid;
	assign forkC_54_out2_ready = brCst_block13_in1_ready;

	assign branchC_56_clk = clk;
	assign branchC_56_rst = rst;
	assign phiC_42_in2_data = branchC_56_out1_data;
	assign phiC_42_in2_valid = branchC_56_out1_valid;
	assign branchC_56_out1_ready = phiC_42_in2_ready;
	assign sink_34_in1_data = branchC_56_out2_data;
	assign sink_34_in1_valid = branchC_56_out2_valid;
	assign branchC_56_out2_ready = sink_34_in1_ready;

	assign source_5_clk = clk;
	assign source_5_rst = rst;
	assign cst_11_in1_data = source_5_out1_data;
	assign cst_11_in1_valid = source_5_out1_valid;
	assign source_5_out1_ready = cst_11_in1_ready;

	assign source_6_clk = clk;
	assign source_6_rst = rst;
	assign cst_12_in1_data = source_6_out1_data;
	assign cst_12_in1_valid = source_6_out1_valid;
	assign source_6_out1_ready = cst_12_in1_ready;

	assign load_43_clk = clk;
	assign load_43_rst = rst;
	assign icmp_44_in1_data = load_43_out1_data;
	assign icmp_44_in1_valid = load_43_out1_valid;
	assign load_43_out1_ready = icmp_44_in1_ready;
	assign MC_pattern_in4_data = load_43_out2_data;
	assign MC_pattern_in4_valid = load_43_out2_valid;
	assign load_43_out2_ready = MC_pattern_in4_ready;

	assign icmp_44_clk = clk;
	assign icmp_44_rst = rst;
	assign fork_36_in1_data = icmp_44_out1_data;
	assign fork_36_in1_valid = icmp_44_out1_valid;
	assign icmp_44_out1_ready = fork_36_in1_ready;

	assign phi_n21_clk = clk;
	assign phi_n21_rst = rst;
	assign fork_20_in1_data = phi_n21_out1_data;
	assign fork_20_in1_valid = phi_n21_out1_valid;
	assign phi_n21_out1_ready = fork_20_in1_ready;

	assign phi_n22_clk = clk;
	assign phi_n22_rst = rst;
	assign fork_21_in1_data = phi_n22_out1_data;
	assign fork_21_in1_valid = phi_n22_out1_valid;
	assign phi_n22_out1_ready = fork_21_in1_ready;

	assign phi_n23_clk = clk;
	assign phi_n23_rst = rst;
	assign branch_29_in1_data = phi_n23_out1_data;
	assign branch_29_in1_valid = phi_n23_out1_valid;
	assign phi_n23_out1_ready = branch_29_in1_ready;

	assign phi_n24_clk = clk;
	assign phi_n24_rst = rst;
	assign branch_30_in1_data = phi_n24_out1_data;
	assign branch_30_in1_valid = phi_n24_out1_valid;
	assign phi_n24_out1_ready = branch_30_in1_ready;

	assign fork_20_clk = clk;
	assign fork_20_rst = rst;
	assign load_43_in2_data = fork_20_out1_data;
	assign load_43_in2_valid = fork_20_out1_valid;
	assign fork_20_out1_ready = load_43_in2_ready;
	assign branch_27_in1_data = fork_20_out2_data;
	assign branch_27_in1_valid = fork_20_out2_valid;
	assign fork_20_out2_ready = branch_27_in1_ready;

	assign fork_21_clk = clk;
	assign fork_21_rst = rst;
	assign icmp_44_in2_data = fork_21_out1_data;
	assign icmp_44_in2_valid = fork_21_out1_valid;
	assign fork_21_out1_ready = icmp_44_in2_ready;
	assign branch_28_in1_data = fork_21_out2_data;
	assign branch_28_in1_valid = fork_21_out2_valid;
	assign fork_21_out2_ready = branch_28_in1_ready;

	assign branch_27_clk = clk;
	assign branch_27_rst = rst;
	assign phi_n25_in2_data = branch_27_out1_data;
	assign phi_n25_in2_valid = branch_27_out1_valid;
	assign branch_27_out1_ready = phi_n25_in2_ready;
	assign phi_n17_in1_data = branch_27_out2_data;
	assign phi_n17_in1_valid = branch_27_out2_valid;
	assign branch_27_out2_ready = phi_n17_in1_ready;

	assign branch_28_clk = clk;
	assign branch_28_rst = rst;
	assign phi_n26_in2_data = branch_28_out1_data;
	assign phi_n26_in2_valid = branch_28_out1_valid;
	assign branch_28_out1_ready = phi_n26_in2_ready;
	assign phi_n18_in1_data = branch_28_out2_data;
	assign phi_n18_in1_valid = branch_28_out2_valid;
	assign branch_28_out2_ready = phi_n18_in1_ready;

	assign branch_29_clk = clk;
	assign branch_29_rst = rst;
	assign phi_n27_in2_data = branch_29_out1_data;
	assign phi_n27_in2_valid = branch_29_out1_valid;
	assign branch_29_out1_ready = phi_n27_in2_ready;
	assign phi_n19_in1_data = branch_29_out2_data;
	assign phi_n19_in1_valid = branch_29_out2_valid;
	assign branch_29_out2_ready = phi_n19_in1_ready;

	assign branch_30_clk = clk;
	assign branch_30_rst = rst;
	assign phi_n28_in2_data = branch_30_out1_data;
	assign phi_n28_in2_valid = branch_30_out1_valid;
	assign branch_30_out1_ready = phi_n28_in2_ready;
	assign phi_n20_in1_data = branch_30_out2_data;
	assign phi_n20_in1_valid = branch_30_out2_valid;
	assign branch_30_out2_ready = phi_n20_in1_ready;

	assign fork_36_clk = clk;
	assign fork_36_rst = rst;
	assign branch_30_in2_data = fork_36_out1_data;
	assign branch_30_in2_valid = fork_36_out1_valid;
	assign fork_36_out1_ready = branch_30_in2_ready;
	assign branch_29_in2_data = fork_36_out2_data;
	assign branch_29_in2_valid = fork_36_out2_valid;
	assign fork_36_out2_ready = branch_29_in2_ready;
	assign branch_28_in2_data = fork_36_out3_data;
	assign branch_28_in2_valid = fork_36_out3_valid;
	assign fork_36_out3_ready = branch_28_in2_ready;
	assign branch_27_in2_data = fork_36_out4_data;
	assign branch_27_in2_valid = fork_36_out4_valid;
	assign fork_36_out4_ready = branch_27_in2_ready;
	assign branchC_53_in2_data = fork_36_out5_data;
	assign branchC_53_in2_valid = fork_36_out5_valid;
	assign fork_36_out5_ready = branchC_53_in2_ready;

	assign phiC_38_clk = clk;
	assign phiC_38_rst = rst;
	assign branchC_53_in1_data = phiC_38_out1_data;
	assign branchC_53_in1_valid = phiC_38_out1_valid;
	assign phiC_38_out1_ready = branchC_53_in1_ready;

	assign branchC_53_clk = clk;
	assign branchC_53_rst = rst;
	assign phiC_40_in2_data = branchC_53_out1_data;
	assign phiC_40_in2_valid = branchC_53_out1_valid;
	assign branchC_53_out1_ready = phiC_40_in2_ready;
	assign phiC_39_in1_data = branchC_53_out2_data;
	assign phiC_39_in1_valid = branchC_53_out2_valid;
	assign branchC_53_out2_ready = phiC_39_in1_ready;

	assign MC_kmpNext_clk = clk;
	assign MC_kmpNext_rst = rst;
	assign kmpNext_ce0 = kmpNext_we0;
	assign load_17_in1_data = MC_kmpNext_out1_data;
	assign load_17_in1_valid = MC_kmpNext_out1_valid;
	assign MC_kmpNext_out1_ready = load_17_in1_ready;
	assign load_48_in1_data = MC_kmpNext_out2_data;
	assign load_48_in1_valid = MC_kmpNext_out2_valid;
	assign MC_kmpNext_out2_ready = load_48_in1_ready;
	assign load_62_in1_data = MC_kmpNext_out3_data;
	assign load_62_in1_valid = MC_kmpNext_out3_valid;
	assign MC_kmpNext_out3_ready = load_62_in1_ready;
	assign end_0_in1_data = MC_kmpNext_out4_data;
	assign end_0_in1_valid = MC_kmpNext_out4_valid;
	assign MC_kmpNext_out4_ready = end_0_in1_ready;

	assign MC_pattern_clk = clk;
	assign MC_pattern_rst = rst;
	assign pattern_ce0 = pattern_we0;
	assign MC_pattern_in6_valid = 0;
	assign MC_pattern_in6_data = 0;
	assign load_5_in1_data = MC_pattern_out1_data;
	assign load_5_in1_valid = MC_pattern_out1_valid;
	assign MC_pattern_out1_ready = load_5_in1_ready;
	assign load_12_in1_data = MC_pattern_out2_data;
	assign load_12_in1_valid = MC_pattern_out2_valid;
	assign MC_pattern_out2_ready = load_12_in1_ready;
	assign load_21_in1_data = MC_pattern_out3_data;
	assign load_21_in1_valid = MC_pattern_out3_valid;
	assign MC_pattern_out3_ready = load_21_in1_ready;
	assign load_43_in1_data = MC_pattern_out4_data;
	assign load_43_in1_valid = MC_pattern_out4_valid;
	assign MC_pattern_out4_ready = load_43_in1_ready;
	assign load_52_in1_data = MC_pattern_out5_data;
	assign load_52_in1_valid = MC_pattern_out5_valid;
	assign MC_pattern_out5_ready = load_52_in1_ready;
	assign end_0_in2_data = MC_pattern_out6_data;
	assign end_0_in2_valid = MC_pattern_out6_valid;
	assign MC_pattern_out6_ready = end_0_in2_ready;

	assign MC_input_clk = clk;
	assign MC_input_rst = rst;
	assign input_ce0 = input_we0;
	assign MC_input_in2_valid = 0;
	assign MC_input_in2_data = 0;
	assign load_36_in1_data = MC_input_out1_data;
	assign load_36_in1_valid = MC_input_out1_valid;
	assign MC_input_out1_ready = load_36_in1_ready;
	assign end_0_in3_data = MC_input_out2_data;
	assign end_0_in3_valid = MC_input_out2_valid;
	assign MC_input_out2_ready = end_0_in3_ready;

	assign sink_1_clk = clk;
	assign sink_1_rst = rst;

	assign sink_2_clk = clk;
	assign sink_2_rst = rst;

	assign sink_3_clk = clk;
	assign sink_3_rst = rst;

	assign sink_4_clk = clk;
	assign sink_4_rst = rst;

	assign sink_5_clk = clk;
	assign sink_5_rst = rst;

	assign sink_6_clk = clk;
	assign sink_6_rst = rst;

	assign sink_7_clk = clk;
	assign sink_7_rst = rst;

	assign sink_8_clk = clk;
	assign sink_8_rst = rst;

	assign sink_9_clk = clk;
	assign sink_9_rst = rst;

	assign sink_10_clk = clk;
	assign sink_10_rst = rst;

	assign sink_11_clk = clk;
	assign sink_11_rst = rst;

	assign sink_12_clk = clk;
	assign sink_12_rst = rst;

	assign sink_13_clk = clk;
	assign sink_13_rst = rst;

	assign sink_14_clk = clk;
	assign sink_14_rst = rst;

	assign sink_15_clk = clk;
	assign sink_15_rst = rst;

	assign sink_16_clk = clk;
	assign sink_16_rst = rst;

	assign sink_17_clk = clk;
	assign sink_17_rst = rst;

	assign sink_18_clk = clk;
	assign sink_18_rst = rst;

	assign sink_19_clk = clk;
	assign sink_19_rst = rst;

	assign sink_20_clk = clk;
	assign sink_20_rst = rst;

	assign sink_21_clk = clk;
	assign sink_21_rst = rst;

	assign sink_22_clk = clk;
	assign sink_22_rst = rst;

	assign sink_23_clk = clk;
	assign sink_23_rst = rst;

	assign sink_24_clk = clk;
	assign sink_24_rst = rst;

	assign sink_25_clk = clk;
	assign sink_25_rst = rst;

	assign sink_26_clk = clk;
	assign sink_26_rst = rst;

	assign sink_27_clk = clk;
	assign sink_27_rst = rst;

	assign sink_28_clk = clk;
	assign sink_28_rst = rst;

	assign sink_29_clk = clk;
	assign sink_29_rst = rst;

	assign sink_30_clk = clk;
	assign sink_30_rst = rst;

	assign sink_31_clk = clk;
	assign sink_31_rst = rst;

	assign sink_32_clk = clk;
	assign sink_32_rst = rst;

	assign sink_33_clk = clk;
	assign sink_33_rst = rst;

	assign sink_34_clk = clk;
	assign sink_34_rst = rst;

	assign Buffer_100_clk = clk;
	assign Buffer_100_rst = rst;
	assign phi_7_in3_data = Buffer_100_out1_data;
	assign phi_7_in3_valid = Buffer_100_out1_valid;
	assign Buffer_100_out1_ready = phi_7_in3_ready;

	assign Buffer_101_clk = clk;
	assign Buffer_101_rst = rst;
	assign phi_n6_in2_data = Buffer_101_out1_data;
	assign phi_n6_in2_valid = Buffer_101_out1_valid;
	assign Buffer_101_out1_ready = phi_n6_in2_ready;

	assign Buffer_102_clk = clk;
	assign Buffer_102_rst = rst;
	assign phi_n7_in2_data = Buffer_102_out1_data;
	assign phi_n7_in2_valid = Buffer_102_out1_valid;
	assign Buffer_102_out1_ready = phi_n7_in2_ready;

	assign Buffer_103_clk = clk;
	assign Buffer_103_rst = rst;
	assign phiC_31_in2_data = Buffer_103_out1_data;
	assign phiC_31_in2_valid = Buffer_103_out1_valid;
	assign Buffer_103_out1_ready = phiC_31_in2_ready;

	assign Buffer_104_clk = clk;
	assign Buffer_104_rst = rst;
	assign phi_1_in3_data = Buffer_104_out1_data;
	assign phi_1_in3_valid = Buffer_104_out1_valid;
	assign Buffer_104_out1_ready = phi_1_in3_ready;

	assign Buffer_105_clk = clk;
	assign Buffer_105_rst = rst;
	assign phi_2_in3_data = Buffer_105_out1_data;
	assign phi_2_in3_valid = Buffer_105_out1_valid;
	assign Buffer_105_out1_ready = phi_2_in3_ready;

	assign Buffer_106_clk = clk;
	assign Buffer_106_rst = rst;
	assign phiC_30_in2_data = Buffer_106_out1_data;
	assign phiC_30_in2_valid = Buffer_106_out1_valid;
	assign Buffer_106_out1_ready = phiC_30_in2_ready;

	assign Buffer_107_clk = clk;
	assign Buffer_107_rst = rst;
	assign phi_38_in3_data = Buffer_107_out1_data;
	assign phi_38_in3_valid = Buffer_107_out1_valid;
	assign Buffer_107_out1_ready = phi_38_in3_ready;

	assign Buffer_108_clk = clk;
	assign Buffer_108_rst = rst;
	assign phi_n10_in2_data = Buffer_108_out1_data;
	assign phi_n10_in2_valid = Buffer_108_out1_valid;
	assign Buffer_108_out1_ready = phi_n10_in2_ready;

	assign Buffer_109_clk = clk;
	assign Buffer_109_rst = rst;
	assign phi_n11_in2_data = Buffer_109_out1_data;
	assign phi_n11_in2_valid = Buffer_109_out1_valid;
	assign Buffer_109_out1_ready = phi_n11_in2_ready;

	assign Buffer_110_clk = clk;
	assign Buffer_110_rst = rst;
	assign phi_n12_in2_data = Buffer_110_out1_data;
	assign phi_n12_in2_valid = Buffer_110_out1_valid;
	assign Buffer_110_out1_ready = phi_n12_in2_ready;

	assign Buffer_111_clk = clk;
	assign Buffer_111_rst = rst;
	assign phiC_37_in2_data = Buffer_111_out1_data;
	assign phiC_37_in2_valid = Buffer_111_out1_valid;
	assign Buffer_111_out1_ready = phiC_37_in2_ready;

	assign Buffer_112_clk = clk;
	assign Buffer_112_rst = rst;
	assign phi_32_in3_data = Buffer_112_out1_data;
	assign phi_32_in3_valid = Buffer_112_out1_valid;
	assign Buffer_112_out1_ready = phi_32_in3_ready;

	assign Buffer_113_clk = clk;
	assign Buffer_113_rst = rst;
	assign phi_31_in3_data = Buffer_113_out1_data;
	assign phi_31_in3_valid = Buffer_113_out1_valid;
	assign Buffer_113_out1_ready = phi_31_in3_ready;

	assign Buffer_114_clk = clk;
	assign Buffer_114_rst = rst;
	assign phi_33_in3_data = Buffer_114_out1_data;
	assign phi_33_in3_valid = Buffer_114_out1_valid;
	assign Buffer_114_out1_ready = phi_33_in3_ready;

	assign Buffer_115_clk = clk;
	assign Buffer_115_rst = rst;
	assign phiC_36_in2_data = Buffer_115_out1_data;
	assign phiC_36_in2_valid = Buffer_115_out1_valid;
	assign Buffer_115_out1_ready = phiC_36_in2_ready;

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_1
		(.clk(phi_1_clk), .rst(phi_1_rst),
		.data_in_bus({{31'b0, phi_1_in1_data}, phi_1_in3_data, phi_1_in2_data}), .valid_in_bus({phi_1_in1_valid, phi_1_in3_valid, phi_1_in2_valid}), .ready_in_bus({phi_1_in1_ready, phi_1_in3_ready, phi_1_in2_ready}), 
		.data_out_bus({phi_1_out1_data}), .valid_out_bus({phi_1_out1_valid}), .ready_out_bus({phi_1_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3), .COND_SIZE(1)) mux_node_phi_2
		(.clk(phi_2_clk), .rst(phi_2_rst),
		.data_in_bus({{2'b0, phi_2_in1_data}, phi_2_in3_data, phi_2_in2_data}), .valid_in_bus({phi_2_in1_valid, phi_2_in3_valid, phi_2_in2_valid}), .ready_in_bus({phi_2_in1_ready, phi_2_in3_ready, phi_2_in2_ready}), 
		.data_out_bus({phi_2_out1_data}), .valid_out_bus({phi_2_out1_valid}), .ready_out_bus({phi_2_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(3), .DATA_SIZE(32)) mc_load_op_load_5
		(.clk(load_5_clk), .rst(load_5_rst),
		.data_in_bus({load_5_in1_data}), .address_in_bus({load_5_in2_data}), .valid_in_bus({load_5_in2_valid, load_5_in1_valid}), .ready_in_bus({load_5_in2_ready, load_5_in1_ready}), 
		.data_out_bus({load_5_out1_data}), .address_out_bus({load_5_out2_data}), .valid_out_bus({load_5_out2_valid, load_5_out1_valid}), .ready_out_bus({load_5_out2_ready, load_5_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block2
		(.clk(brCst_block2_clk), .rst(brCst_block2_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block2_in1_valid}), .ready_in_bus({brCst_block2_in1_ready}), 
		.data_out_bus({brCst_block2_out1_data}), .valid_out_bus({brCst_block2_out1_valid}), .ready_out_bus({brCst_block2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) fork_node_fork_0
		(.clk(fork_0_clk), .rst(fork_0_rst),
		.data_in_bus({fork_0_in1_data}), .valid_in_bus({fork_0_in1_valid}), .ready_in_bus({fork_0_in1_ready}), 
		.data_out_bus({fork_0_out2_data, fork_0_out1_data}), .valid_out_bus({fork_0_out2_valid, fork_0_out1_valid}), .ready_out_bus({fork_0_out2_ready, fork_0_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_2
		(.clk(branch_2_clk), .rst(branch_2_rst),
		.data_in_bus({{31'b0, branch_2_in2_data}, branch_2_in1_data}), .valid_in_bus({branch_2_in2_valid, branch_2_in1_valid}), .ready_in_bus({branch_2_in2_ready, branch_2_in1_ready}), 
		.data_out_bus({branch_2_out2_data, branch_2_out1_data}), .valid_out_bus({branch_2_out2_valid, branch_2_out1_valid}), .ready_out_bus({branch_2_out2_ready, branch_2_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_3
		(.clk(branch_3_clk), .rst(branch_3_rst),
		.data_in_bus({{31'b0, branch_3_in2_data}, branch_3_in1_data}), .valid_in_bus({branch_3_in2_valid, branch_3_in1_valid}), .ready_in_bus({branch_3_in2_ready, branch_3_in1_ready}), 
		.data_out_bus({branch_3_out2_data, branch_3_out1_data}), .valid_out_bus({branch_3_out2_valid, branch_3_out1_valid}), .ready_out_bus({branch_3_out2_ready, branch_3_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) branch_node_branch_4
		(.clk(branch_4_clk), .rst(branch_4_rst),
		.data_in_bus({{2'b0, branch_4_in2_data}, branch_4_in1_data}), .valid_in_bus({branch_4_in2_valid, branch_4_in1_valid}), .ready_in_bus({branch_4_in2_ready, branch_4_in1_ready}), 
		.data_out_bus({branch_4_out2_data, branch_4_out1_data}), .valid_out_bus({branch_4_out2_valid, branch_4_out1_valid}), .ready_out_bus({branch_4_out2_ready, branch_4_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_28
		(.clk(fork_28_clk), .rst(fork_28_rst),
		.data_in_bus({fork_28_in1_data}), .valid_in_bus({fork_28_in1_valid}), .ready_in_bus({fork_28_in1_ready}), 
		.data_out_bus({fork_28_out4_data, fork_28_out3_data, fork_28_out2_data, fork_28_out1_data}), .valid_out_bus({fork_28_out4_valid, fork_28_out3_valid, fork_28_out2_valid, fork_28_out1_valid}), .ready_out_bus({fork_28_out4_ready, fork_28_out3_ready, fork_28_out2_ready, fork_28_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_30
		(.clk(phiC_30_clk), .rst(phiC_30_rst),
		.data_in_bus({phiC_30_in2_data, phiC_30_in1_data}), .valid_in_bus({phiC_30_in2_valid, phiC_30_in1_valid}), .ready_in_bus({phiC_30_in2_ready, phiC_30_in1_ready}), 
		.data_out_bus({phiC_30_out2_data, phiC_30_out1_data}), .valid_out_bus({phiC_30_out2_valid, phiC_30_out1_valid}), .ready_out_bus({phiC_30_out2_ready, phiC_30_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_43
		(.clk(forkC_43_clk), .rst(forkC_43_rst),
		.data_in_bus({forkC_43_in1_data}), .valid_in_bus({forkC_43_in1_valid}), .ready_in_bus({forkC_43_in1_ready}), 
		.data_out_bus({forkC_43_out2_data, forkC_43_out1_data}), .valid_out_bus({forkC_43_out2_valid, forkC_43_out1_valid}), .ready_out_bus({forkC_43_out2_ready, forkC_43_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_45
		(.clk(branchC_45_clk), .rst(branchC_45_rst),
		.data_in_bus({{branchC_45_in2_data}, branchC_45_in1_data}), .valid_in_bus({branchC_45_in2_valid, branchC_45_in1_valid}), .ready_in_bus({branchC_45_in2_ready, branchC_45_in1_ready}), 
		.data_out_bus({branchC_45_out2_data, branchC_45_out1_data}), .valid_out_bus({branchC_45_out2_valid, branchC_45_out1_valid}), .ready_out_bus({branchC_45_out2_ready, branchC_45_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_57
		(.clk(fork_57_clk), .rst(fork_57_rst),
		.data_in_bus({fork_57_in1_data}), .valid_in_bus({fork_57_in1_valid}), .ready_in_bus({fork_57_in1_ready}), 
		.data_out_bus({fork_57_out2_data, fork_57_out1_data}), .valid_out_bus({fork_57_out2_valid, fork_57_out1_valid}), .ready_out_bus({fork_57_out2_ready, fork_57_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_31
		(.clk(phi_31_clk), .rst(phi_31_rst),
		.data_in_bus({{31'b0, phi_31_in1_data}, phi_31_in3_data, phi_31_in2_data}), .valid_in_bus({phi_31_in1_valid, phi_31_in3_valid, phi_31_in2_valid}), .ready_in_bus({phi_31_in1_ready, phi_31_in3_ready, phi_31_in2_ready}), 
		.data_out_bus({phi_31_out1_data}), .valid_out_bus({phi_31_out1_valid}), .ready_out_bus({phi_31_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_32
		(.clk(phi_32_clk), .rst(phi_32_rst),
		.data_in_bus({{31'b0, phi_32_in1_data}, phi_32_in3_data, phi_32_in2_data}), .valid_in_bus({phi_32_in1_valid, phi_32_in3_valid, phi_32_in2_valid}), .ready_in_bus({phi_32_in1_ready, phi_32_in3_ready, phi_32_in2_ready}), 
		.data_out_bus({phi_32_out1_data}), .valid_out_bus({phi_32_out1_valid}), .ready_out_bus({phi_32_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10), .COND_SIZE(1)) mux_node_phi_33
		(.clk(phi_33_clk), .rst(phi_33_rst),
		.data_in_bus({{9'b0, phi_33_in1_data}, phi_33_in3_data, phi_33_in2_data}), .valid_in_bus({phi_33_in1_valid, phi_33_in3_valid, phi_33_in2_valid}), .ready_in_bus({phi_33_in1_ready, phi_33_in3_ready, phi_33_in2_ready}), 
		.data_out_bus({phi_33_out1_data}), .valid_out_bus({phi_33_out1_valid}), .ready_out_bus({phi_33_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(10), .DATA_SIZE(32)) mc_load_op_load_36
		(.clk(load_36_clk), .rst(load_36_rst),
		.data_in_bus({load_36_in1_data}), .address_in_bus({load_36_in2_data}), .valid_in_bus({load_36_in2_valid, load_36_in1_valid}), .ready_in_bus({load_36_in2_ready, load_36_in1_ready}), 
		.data_out_bus({load_36_out1_data}), .address_out_bus({load_36_out2_data}), .valid_out_bus({load_36_out2_valid, load_36_out1_valid}), .ready_out_bus({load_36_out2_ready, load_36_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block8
		(.clk(brCst_block8_clk), .rst(brCst_block8_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block8_in1_valid}), .ready_in_bus({brCst_block8_in1_ready}), 
		.data_out_bus({brCst_block8_out1_data}), .valid_out_bus({brCst_block8_out1_valid}), .ready_out_bus({brCst_block8_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) fork_node_fork_4
		(.clk(fork_4_clk), .rst(fork_4_rst),
		.data_in_bus({fork_4_in1_data}), .valid_in_bus({fork_4_in1_valid}), .ready_in_bus({fork_4_in1_ready}), 
		.data_out_bus({fork_4_out2_data, fork_4_out1_data}), .valid_out_bus({fork_4_out2_valid, fork_4_out1_valid}), .ready_out_bus({fork_4_out2_ready, fork_4_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_19
		(.clk(branch_19_clk), .rst(branch_19_rst),
		.data_in_bus({{31'b0, branch_19_in2_data}, branch_19_in1_data}), .valid_in_bus({branch_19_in2_valid, branch_19_in1_valid}), .ready_in_bus({branch_19_in2_ready, branch_19_in1_ready}), 
		.data_out_bus({branch_19_out2_data, branch_19_out1_data}), .valid_out_bus({branch_19_out2_valid, branch_19_out1_valid}), .ready_out_bus({branch_19_out2_ready, branch_19_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_20
		(.clk(branch_20_clk), .rst(branch_20_rst),
		.data_in_bus({{31'b0, branch_20_in2_data}, branch_20_in1_data}), .valid_in_bus({branch_20_in2_valid, branch_20_in1_valid}), .ready_in_bus({branch_20_in2_ready, branch_20_in1_ready}), 
		.data_out_bus({branch_20_out2_data, branch_20_out1_data}), .valid_out_bus({branch_20_out2_valid, branch_20_out1_valid}), .ready_out_bus({branch_20_out2_ready, branch_20_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_21
		(.clk(branch_21_clk), .rst(branch_21_rst),
		.data_in_bus({{31'b0, branch_21_in2_data}, branch_21_in1_data}), .valid_in_bus({branch_21_in2_valid, branch_21_in1_valid}), .ready_in_bus({branch_21_in2_ready, branch_21_in1_ready}), 
		.data_out_bus({branch_21_out2_data, branch_21_out1_data}), .valid_out_bus({branch_21_out2_valid, branch_21_out1_valid}), .ready_out_bus({branch_21_out2_ready, branch_21_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) branch_node_branch_22
		(.clk(branch_22_clk), .rst(branch_22_rst),
		.data_in_bus({{9'b0, branch_22_in2_data}, branch_22_in1_data}), .valid_in_bus({branch_22_in2_valid, branch_22_in1_valid}), .ready_in_bus({branch_22_in2_ready, branch_22_in1_ready}), 
		.data_out_bus({branch_22_out2_data, branch_22_out1_data}), .valid_out_bus({branch_22_out2_valid, branch_22_out1_valid}), .ready_out_bus({branch_22_out2_ready, branch_22_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_34
		(.clk(fork_34_clk), .rst(fork_34_rst),
		.data_in_bus({fork_34_in1_data}), .valid_in_bus({fork_34_in1_valid}), .ready_in_bus({fork_34_in1_ready}), 
		.data_out_bus({fork_34_out5_data, fork_34_out4_data, fork_34_out3_data, fork_34_out2_data, fork_34_out1_data}), .valid_out_bus({fork_34_out5_valid, fork_34_out4_valid, fork_34_out3_valid, fork_34_out2_valid, fork_34_out1_valid}), .ready_out_bus({fork_34_out5_ready, fork_34_out4_ready, fork_34_out3_ready, fork_34_out2_ready, fork_34_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_36
		(.clk(phiC_36_clk), .rst(phiC_36_rst),
		.data_in_bus({phiC_36_in2_data, phiC_36_in1_data}), .valid_in_bus({phiC_36_in2_valid, phiC_36_in1_valid}), .ready_in_bus({phiC_36_in2_ready, phiC_36_in1_ready}), 
		.data_out_bus({phiC_36_out2_data, phiC_36_out1_data}), .valid_out_bus({phiC_36_out2_valid, phiC_36_out1_valid}), .ready_out_bus({phiC_36_out2_ready, phiC_36_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_49
		(.clk(forkC_49_clk), .rst(forkC_49_rst),
		.data_in_bus({forkC_49_in1_data}), .valid_in_bus({forkC_49_in1_valid}), .ready_in_bus({forkC_49_in1_ready}), 
		.data_out_bus({forkC_49_out2_data, forkC_49_out1_data}), .valid_out_bus({forkC_49_out2_valid, forkC_49_out1_valid}), .ready_out_bus({forkC_49_out2_ready, forkC_49_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_51
		(.clk(branchC_51_clk), .rst(branchC_51_rst),
		.data_in_bus({{branchC_51_in2_data}, branchC_51_in1_data}), .valid_in_bus({branchC_51_in2_valid, branchC_51_in1_valid}), .ready_in_bus({branchC_51_in2_ready, branchC_51_in1_ready}), 
		.data_out_bus({branchC_51_out2_data, branchC_51_out1_data}), .valid_out_bus({branchC_51_out2_valid, branchC_51_out1_valid}), .ready_out_bus({branchC_51_out2_ready, branchC_51_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_59
		(.clk(fork_59_clk), .rst(fork_59_rst),
		.data_in_bus({fork_59_in1_data}), .valid_in_bus({fork_59_in1_valid}), .ready_in_bus({fork_59_in1_ready}), 
		.data_out_bus({fork_59_out3_data, fork_59_out2_data, fork_59_out1_data}), .valid_out_bus({fork_59_out3_valid, fork_59_out2_valid, fork_59_out1_valid}), .ready_out_bus({fork_59_out3_ready, fork_59_out2_ready, fork_59_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(32), .DATA_SIZE(32)) mc_load_op_load_48
		(.clk(load_48_clk), .rst(load_48_rst),
		.data_in_bus({load_48_in1_data}), .address_in_bus({load_48_in2_data}), .valid_in_bus({load_48_in2_valid, load_48_in1_valid}), .ready_in_bus({load_48_in2_ready, load_48_in1_ready}), 
		.data_out_bus({load_48_out1_data}), .address_out_bus({load_48_out2_data}), .valid_out_bus({load_48_out2_valid, load_48_out1_valid}), .ready_out_bus({load_48_out2_ready, load_48_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block11
		(.clk(brCst_block11_clk), .rst(brCst_block11_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block11_in1_valid}), .ready_in_bus({brCst_block11_in1_ready}), 
		.data_out_bus({brCst_block11_out1_data}), .valid_out_bus({brCst_block11_out1_valid}), .ready_out_bus({brCst_block11_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n17
		(.clk(phi_n17_clk), .rst(phi_n17_rst),
		.data_in_bus({phi_n17_in1_data}), .valid_in_bus({phi_n17_in1_valid}), .ready_in_bus({phi_n17_in1_ready}), 
		.data_out_bus({phi_n17_out1_data}), .valid_out_bus({phi_n17_out1_valid}), .ready_out_bus({phi_n17_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n18
		(.clk(phi_n18_clk), .rst(phi_n18_rst),
		.data_in_bus({phi_n18_in1_data}), .valid_in_bus({phi_n18_in1_valid}), .ready_in_bus({phi_n18_in1_ready}), 
		.data_out_bus({phi_n18_out1_data}), .valid_out_bus({phi_n18_out1_valid}), .ready_out_bus({phi_n18_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n19
		(.clk(phi_n19_clk), .rst(phi_n19_rst),
		.data_in_bus({phi_n19_in1_data}), .valid_in_bus({phi_n19_in1_valid}), .ready_in_bus({phi_n19_in1_ready}), 
		.data_out_bus({phi_n19_out1_data}), .valid_out_bus({phi_n19_out1_valid}), .ready_out_bus({phi_n19_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) merge_node_phi_n20
		(.clk(phi_n20_clk), .rst(phi_n20_rst),
		.data_in_bus({phi_n20_in1_data}), .valid_in_bus({phi_n20_in1_valid}), .ready_in_bus({phi_n20_in1_ready}), 
		.data_out_bus({phi_n20_out1_data}), .valid_out_bus({phi_n20_out1_valid}), .ready_out_bus({phi_n20_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_31
		(.clk(branch_31_clk), .rst(branch_31_rst),
		.data_in_bus({{31'b0, branch_31_in2_data}, branch_31_in1_data}), .valid_in_bus({branch_31_in2_valid, branch_31_in1_valid}), .ready_in_bus({branch_31_in2_ready, branch_31_in1_ready}), 
		.data_out_bus({branch_31_out2_data, branch_31_out1_data}), .valid_out_bus({branch_31_out2_valid, branch_31_out1_valid}), .ready_out_bus({branch_31_out2_ready, branch_31_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_32
		(.clk(branch_32_clk), .rst(branch_32_rst),
		.data_in_bus({{31'b0, branch_32_in2_data}, branch_32_in1_data}), .valid_in_bus({branch_32_in2_valid, branch_32_in1_valid}), .ready_in_bus({branch_32_in2_ready, branch_32_in1_ready}), 
		.data_out_bus({branch_32_out2_data, branch_32_out1_data}), .valid_out_bus({branch_32_out2_valid, branch_32_out1_valid}), .ready_out_bus({branch_32_out2_ready, branch_32_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_33
		(.clk(branch_33_clk), .rst(branch_33_rst),
		.data_in_bus({{31'b0, branch_33_in2_data}, branch_33_in1_data}), .valid_in_bus({branch_33_in2_valid, branch_33_in1_valid}), .ready_in_bus({branch_33_in2_ready, branch_33_in1_ready}), 
		.data_out_bus({branch_33_out2_data, branch_33_out1_data}), .valid_out_bus({branch_33_out2_valid, branch_33_out1_valid}), .ready_out_bus({branch_33_out2_ready, branch_33_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) branch_node_branch_34
		(.clk(branch_34_clk), .rst(branch_34_rst),
		.data_in_bus({{9'b0, branch_34_in2_data}, branch_34_in1_data}), .valid_in_bus({branch_34_in2_valid, branch_34_in1_valid}), .ready_in_bus({branch_34_in2_ready, branch_34_in1_ready}), 
		.data_out_bus({branch_34_out2_data, branch_34_out1_data}), .valid_out_bus({branch_34_out2_valid, branch_34_out1_valid}), .ready_out_bus({branch_34_out2_ready, branch_34_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_37
		(.clk(fork_37_clk), .rst(fork_37_rst),
		.data_in_bus({fork_37_in1_data}), .valid_in_bus({fork_37_in1_valid}), .ready_in_bus({fork_37_in1_ready}), 
		.data_out_bus({fork_37_out5_data, fork_37_out4_data, fork_37_out3_data, fork_37_out2_data, fork_37_out1_data}), .valid_out_bus({fork_37_out5_valid, fork_37_out4_valid, fork_37_out3_valid, fork_37_out2_valid, fork_37_out1_valid}), .ready_out_bus({fork_37_out5_ready, fork_37_out4_ready, fork_37_out3_ready, fork_37_out2_ready, fork_37_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_39
		(.clk(phiC_39_clk), .rst(phiC_39_rst),
		.data_in_bus({phiC_39_in1_data}), .valid_in_bus({phiC_39_in1_valid}), .ready_in_bus({phiC_39_in1_ready}), 
		.data_out_bus({phiC_39_out1_data}), .valid_out_bus({phiC_39_out1_valid}), .ready_out_bus({phiC_39_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_52
		(.clk(forkC_52_clk), .rst(forkC_52_rst),
		.data_in_bus({forkC_52_in1_data}), .valid_in_bus({forkC_52_in1_valid}), .ready_in_bus({forkC_52_in1_ready}), 
		.data_out_bus({forkC_52_out2_data, forkC_52_out1_data}), .valid_out_bus({forkC_52_out2_valid, forkC_52_out1_valid}), .ready_out_bus({forkC_52_out2_ready, forkC_52_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_54
		(.clk(branchC_54_clk), .rst(branchC_54_rst),
		.data_in_bus({{branchC_54_in2_data}, branchC_54_in1_data}), .valid_in_bus({branchC_54_in2_valid, branchC_54_in1_valid}), .ready_in_bus({branchC_54_in2_ready, branchC_54_in1_ready}), 
		.data_out_bus({branchC_54_out2_data, branchC_54_out1_data}), .valid_out_bus({branchC_54_out2_valid, branchC_54_out1_valid}), .ready_out_bus({branchC_54_out2_ready, branchC_54_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(32), .DATA_SIZE(32)) mc_load_op_load_52
		(.clk(load_52_clk), .rst(load_52_rst),
		.data_in_bus({load_52_in1_data}), .address_in_bus({load_52_in2_data}), .valid_in_bus({load_52_in2_valid, load_52_in1_valid}), .ready_in_bus({load_52_in2_ready, load_52_in1_ready}), 
		.data_out_bus({load_52_out1_data}), .address_out_bus({load_52_out2_data}), .valid_out_bus({load_52_out2_valid, load_52_out1_valid}), .ready_out_bus({load_52_out2_ready, load_52_out1_ready}));

	icmp_eq_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(1)) icmp_eq_op_icmp_53
		(.clk(icmp_53_clk), .rst(icmp_53_rst),
		.data_in_bus({icmp_53_in2_data, icmp_53_in1_data}), .valid_in_bus({icmp_53_in2_valid, icmp_53_in1_valid}), .ready_in_bus({icmp_53_in2_ready, icmp_53_in1_ready}), 
		.data_out_bus({icmp_53_out1_data}), .valid_out_bus({icmp_53_out1_valid}), .ready_out_bus({icmp_53_out1_ready}));

	zext_op #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) zext_op_zext_54
		(.clk(zext_54_clk), .rst(zext_54_rst),
		.data_in_bus({zext_54_in1_data}), .valid_in_bus({zext_54_in1_valid}), .ready_in_bus({zext_54_in1_ready}), 
		.data_out_bus({zext_54_out1_data}), .valid_out_bus({zext_54_out1_valid}), .ready_out_bus({zext_54_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_55
		(.clk(add_55_clk), .rst(add_55_rst),
		.data_in_bus({add_55_in2_data, add_55_in1_data}), .valid_in_bus({add_55_in2_valid, add_55_in1_valid}), .ready_in_bus({add_55_in2_ready, add_55_in1_ready}), 
		.data_out_bus({add_55_out1_data}), .valid_out_bus({add_55_out1_valid}), .ready_out_bus({add_55_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(2), .DATA_OUT_SIZE(2)) const_node_cst_10
		(.clk(cst_10_clk), .rst(cst_10_rst),
		.data_in_bus({2'd3}), .valid_in_bus({cst_10_in1_valid}), .ready_in_bus({cst_10_in1_ready}), 
		.data_out_bus({cst_10_out1_data}), .valid_out_bus({cst_10_out1_valid}), .ready_out_bus({cst_10_out1_ready}));

	icmp_sgt_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(1)) icmp_sgt_op_icmp_56
		(.clk(icmp_56_clk), .rst(icmp_56_rst),
		.data_in_bus({icmp_56_in2_data, icmp_56_in1_data}), .valid_in_bus({icmp_56_in2_valid, icmp_56_in1_valid}), .ready_in_bus({icmp_56_in2_ready, icmp_56_in1_ready}), 
		.data_out_bus({icmp_56_out1_data}), .valid_out_bus({icmp_56_out1_valid}), .ready_out_bus({icmp_56_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n25
		(.clk(phi_n25_clk), .rst(phi_n25_rst),
		.data_in_bus({phi_n25_in2_data, phi_n25_in1_data}), .valid_in_bus({phi_n25_in2_valid, phi_n25_in1_valid}), .ready_in_bus({phi_n25_in2_ready, phi_n25_in1_ready}), 
		.data_out_bus({phi_n25_out1_data}), .valid_out_bus({phi_n25_out1_valid}), .ready_out_bus({phi_n25_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n26
		(.clk(phi_n26_clk), .rst(phi_n26_rst),
		.data_in_bus({phi_n26_in2_data, phi_n26_in1_data}), .valid_in_bus({phi_n26_in2_valid, phi_n26_in1_valid}), .ready_in_bus({phi_n26_in2_ready, phi_n26_in1_ready}), 
		.data_out_bus({phi_n26_out1_data}), .valid_out_bus({phi_n26_out1_valid}), .ready_out_bus({phi_n26_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n27
		(.clk(phi_n27_clk), .rst(phi_n27_rst),
		.data_in_bus({phi_n27_in2_data, phi_n27_in1_data}), .valid_in_bus({phi_n27_in2_valid, phi_n27_in1_valid}), .ready_in_bus({phi_n27_in2_ready, phi_n27_in1_ready}), 
		.data_out_bus({phi_n27_out1_data}), .valid_out_bus({phi_n27_out1_valid}), .ready_out_bus({phi_n27_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) merge_node_phi_n28
		(.clk(phi_n28_clk), .rst(phi_n28_rst),
		.data_in_bus({phi_n28_in2_data, phi_n28_in1_data}), .valid_in_bus({phi_n28_in2_valid, phi_n28_in1_valid}), .ready_in_bus({phi_n28_in2_ready, phi_n28_in1_ready}), 
		.data_out_bus({phi_n28_out1_data}), .valid_out_bus({phi_n28_out1_valid}), .ready_out_bus({phi_n28_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_6
		(.clk(fork_6_clk), .rst(fork_6_rst),
		.data_in_bus({fork_6_in1_data}), .valid_in_bus({fork_6_in1_valid}), .ready_in_bus({fork_6_in1_ready}), 
		.data_out_bus({fork_6_out2_data, fork_6_out1_data}), .valid_out_bus({fork_6_out2_valid, fork_6_out1_valid}), .ready_out_bus({fork_6_out2_ready, fork_6_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_24
		(.clk(fork_24_clk), .rst(fork_24_rst),
		.data_in_bus({fork_24_in1_data}), .valid_in_bus({fork_24_in1_valid}), .ready_in_bus({fork_24_in1_ready}), 
		.data_out_bus({fork_24_out2_data, fork_24_out1_data}), .valid_out_bus({fork_24_out2_valid, fork_24_out1_valid}), .ready_out_bus({fork_24_out2_ready, fork_24_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_35
		(.clk(branch_35_clk), .rst(branch_35_rst),
		.data_in_bus({{31'b0, branch_35_in2_data}, branch_35_in1_data}), .valid_in_bus({branch_35_in2_valid, branch_35_in1_valid}), .ready_in_bus({branch_35_in2_ready, branch_35_in1_ready}), 
		.data_out_bus({branch_35_out2_data, branch_35_out1_data}), .valid_out_bus({branch_35_out2_valid, branch_35_out1_valid}), .ready_out_bus({branch_35_out2_ready, branch_35_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_36
		(.clk(branch_36_clk), .rst(branch_36_rst),
		.data_in_bus({{31'b0, branch_36_in2_data}, branch_36_in1_data}), .valid_in_bus({branch_36_in2_valid, branch_36_in1_valid}), .ready_in_bus({branch_36_in2_ready, branch_36_in1_ready}), 
		.data_out_bus({branch_36_out2_data, branch_36_out1_data}), .valid_out_bus({branch_36_out2_valid, branch_36_out1_valid}), .ready_out_bus({branch_36_out2_ready, branch_36_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) branch_node_branch_37
		(.clk(branch_37_clk), .rst(branch_37_rst),
		.data_in_bus({{9'b0, branch_37_in2_data}, branch_37_in1_data}), .valid_in_bus({branch_37_in2_valid, branch_37_in1_valid}), .ready_in_bus({branch_37_in2_ready, branch_37_in1_ready}), 
		.data_out_bus({branch_37_out2_data, branch_37_out1_data}), .valid_out_bus({branch_37_out2_valid, branch_37_out1_valid}), .ready_out_bus({branch_37_out2_ready, branch_37_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_38
		(.clk(fork_38_clk), .rst(fork_38_rst),
		.data_in_bus({fork_38_in1_data}), .valid_in_bus({fork_38_in1_valid}), .ready_in_bus({fork_38_in1_ready}), 
		.data_out_bus({fork_38_out4_data, fork_38_out3_data, fork_38_out2_data, fork_38_out1_data}), .valid_out_bus({fork_38_out4_valid, fork_38_out3_valid, fork_38_out2_valid, fork_38_out1_valid}), .ready_out_bus({fork_38_out4_ready, fork_38_out3_ready, fork_38_out2_ready, fork_38_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_40
		(.clk(phiC_40_clk), .rst(phiC_40_rst),
		.data_in_bus({phiC_40_in2_data, phiC_40_in1_data}), .valid_in_bus({phiC_40_in2_valid, phiC_40_in1_valid}), .ready_in_bus({phiC_40_in2_ready, phiC_40_in1_ready}), 
		.data_out_bus({phiC_40_out1_data}), .valid_out_bus({phiC_40_out1_valid}), .ready_out_bus({phiC_40_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_55
		(.clk(branchC_55_clk), .rst(branchC_55_rst),
		.data_in_bus({{branchC_55_in2_data}, branchC_55_in1_data}), .valid_in_bus({branchC_55_in2_valid, branchC_55_in1_valid}), .ready_in_bus({branchC_55_in2_ready, branchC_55_in1_ready}), 
		.data_out_bus({branchC_55_out2_data, branchC_55_out1_data}), .valid_out_bus({branchC_55_out2_valid, branchC_55_out1_valid}), .ready_out_bus({branchC_55_out2_ready, branchC_55_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(2))source_node_source_4
		(.clk(source_4_clk), .rst(source_4_rst),
		.data_out_bus({source_4_out1_data}), .valid_out_bus({source_4_out1_valid}), .ready_out_bus({source_4_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_0
		(.clk(cst_0_clk), .rst(cst_0_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_0_in1_valid}), .ready_in_bus({cst_0_in1_ready}), 
		.data_out_bus({cst_0_out1_data}), .valid_out_bus({cst_0_out1_valid}), .ready_out_bus({cst_0_out1_ready}));

	mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(1), .DATA_SIZE(1)) mc_store_op_store_0
		(.clk(store_0_clk), .rst(store_0_rst),
		.data_in_bus({store_0_in1_data}), .address_in_bus({store_0_in2_data}), .valid_in_bus({store_0_in2_valid, store_0_in1_valid}), .ready_in_bus({store_0_in2_ready, store_0_in1_ready}), 
		.data_out_bus({store_0_out1_data}), .address_out_bus({store_0_out2_data}), .valid_out_bus({store_0_out2_valid, store_0_out1_valid}), .ready_out_bus({store_0_out2_ready, store_0_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block1
		(.clk(brCst_block1_clk), .rst(brCst_block1_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block1_in1_valid}), .ready_in_bus({brCst_block1_in1_ready}), 
		.data_out_bus({brCst_block1_out1_data}), .valid_out_bus({brCst_block1_out1_valid}), .ready_out_bus({brCst_block1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_1
		(.clk(cst_1_clk), .rst(cst_1_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_1_in1_valid}), .ready_in_bus({cst_1_in1_ready}), 
		.data_out_bus({cst_1_out1_data}), .valid_out_bus({cst_1_out1_valid}), .ready_out_bus({cst_1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_2
		(.clk(cst_2_clk), .rst(cst_2_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_2_in1_valid}), .ready_in_bus({cst_2_in1_ready}), 
		.data_out_bus({cst_2_out1_data}), .valid_out_bus({cst_2_out1_valid}), .ready_out_bus({cst_2_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_15
		(.clk(cst_15_clk), .rst(cst_15_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_15_in1_valid}), .ready_in_bus({cst_15_in1_ready}), 
		.data_out_bus({cst_15_out1_data}), .valid_out_bus({cst_15_out1_valid}), .ready_out_bus({cst_15_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_0
		(.clk(branch_0_clk), .rst(branch_0_rst),
		.data_in_bus({{branch_0_in2_data}, branch_0_in1_data}), .valid_in_bus({branch_0_in2_valid, branch_0_in1_valid}), .ready_in_bus({branch_0_in2_ready, branch_0_in1_ready}), 
		.data_out_bus({branch_0_out2_data, branch_0_out1_data}), .valid_out_bus({branch_0_out2_valid, branch_0_out1_valid}), .ready_out_bus({branch_0_out2_ready, branch_0_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_1
		(.clk(branch_1_clk), .rst(branch_1_rst),
		.data_in_bus({{branch_1_in2_data}, branch_1_in1_data}), .valid_in_bus({branch_1_in2_valid, branch_1_in1_valid}), .ready_in_bus({branch_1_in2_ready, branch_1_in1_ready}), 
		.data_out_bus({branch_1_out2_data, branch_1_out1_data}), .valid_out_bus({branch_1_out2_valid, branch_1_out1_valid}), .ready_out_bus({branch_1_out2_ready, branch_1_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_27
		(.clk(fork_27_clk), .rst(fork_27_rst),
		.data_in_bus({fork_27_in1_data}), .valid_in_bus({fork_27_in1_valid}), .ready_in_bus({fork_27_in1_ready}), 
		.data_out_bus({fork_27_out3_data, fork_27_out2_data, fork_27_out1_data}), .valid_out_bus({fork_27_out3_valid, fork_27_out2_valid, fork_27_out1_valid}), .ready_out_bus({fork_27_out3_ready, fork_27_out2_ready, fork_27_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_16
		(.clk(cst_16_clk), .rst(cst_16_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_16_in1_valid}), .ready_in_bus({cst_16_in1_ready}), 
		.data_out_bus({cst_16_out1_data}), .valid_out_bus({cst_16_out1_valid}), .ready_out_bus({cst_16_out1_ready}));

	start_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) start_node_start_0
		(.clk(start_0_clk), .rst(start_0_rst),
		.data_in_bus({start_0_in1_data}), .valid_in_bus({start_0_in1_valid}), .ready_in_bus({start_0_in1_ready}), 
		.data_out_bus({start_0_out1_data}), .valid_out_bus({start_0_out1_valid}), .ready_out_bus({start_0_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(7), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_42
		(.clk(forkC_42_clk), .rst(forkC_42_rst),
		.data_in_bus({forkC_42_in1_data}), .valid_in_bus({forkC_42_in1_valid}), .ready_in_bus({forkC_42_in1_ready}), 
		.data_out_bus({forkC_42_out7_data, forkC_42_out6_data, forkC_42_out5_data, forkC_42_out4_data, forkC_42_out3_data, forkC_42_out2_data, forkC_42_out1_data}), .valid_out_bus({forkC_42_out7_valid, forkC_42_out6_valid, forkC_42_out5_valid, forkC_42_out4_valid, forkC_42_out3_valid, forkC_42_out2_valid, forkC_42_out1_valid}), .ready_out_bus({forkC_42_out7_ready, forkC_42_out6_ready, forkC_42_out5_ready, forkC_42_out4_ready, forkC_42_out3_ready, forkC_42_out2_ready, forkC_42_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_44
		(.clk(branchC_44_clk), .rst(branchC_44_rst),
		.data_in_bus({{branchC_44_in2_data}, branchC_44_in1_data}), .valid_in_bus({branchC_44_in2_valid, branchC_44_in1_valid}), .ready_in_bus({branchC_44_in2_ready, branchC_44_in1_ready}), 
		.data_out_bus({branchC_44_out2_data, branchC_44_out1_data}), .valid_out_bus({branchC_44_out2_valid, branchC_44_out1_valid}), .ready_out_bus({branchC_44_out2_ready, branchC_44_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block7
		(.clk(brCst_block7_clk), .rst(brCst_block7_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block7_in1_valid}), .ready_in_bus({brCst_block7_in1_ready}), 
		.data_out_bus({brCst_block7_out1_data}), .valid_out_bus({brCst_block7_out1_valid}), .ready_out_bus({brCst_block7_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_6
		(.clk(cst_6_clk), .rst(cst_6_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_6_in1_valid}), .ready_in_bus({cst_6_in1_ready}), 
		.data_out_bus({cst_6_out1_data}), .valid_out_bus({cst_6_out1_valid}), .ready_out_bus({cst_6_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_7
		(.clk(cst_7_clk), .rst(cst_7_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_7_in1_valid}), .ready_in_bus({cst_7_in1_ready}), 
		.data_out_bus({cst_7_out1_data}), .valid_out_bus({cst_7_out1_valid}), .ready_out_bus({cst_7_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_8
		(.clk(cst_8_clk), .rst(cst_8_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_8_in1_valid}), .ready_in_bus({cst_8_in1_ready}), 
		.data_out_bus({cst_8_out1_data}), .valid_out_bus({cst_8_out1_valid}), .ready_out_bus({cst_8_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_16
		(.clk(branch_16_clk), .rst(branch_16_rst),
		.data_in_bus({{branch_16_in2_data}, branch_16_in1_data}), .valid_in_bus({branch_16_in2_valid, branch_16_in1_valid}), .ready_in_bus({branch_16_in2_ready, branch_16_in1_ready}), 
		.data_out_bus({branch_16_out2_data, branch_16_out1_data}), .valid_out_bus({branch_16_out2_valid, branch_16_out1_valid}), .ready_out_bus({branch_16_out2_ready, branch_16_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_17
		(.clk(branch_17_clk), .rst(branch_17_rst),
		.data_in_bus({{branch_17_in2_data}, branch_17_in1_data}), .valid_in_bus({branch_17_in2_valid, branch_17_in1_valid}), .ready_in_bus({branch_17_in2_ready, branch_17_in1_ready}), 
		.data_out_bus({branch_17_out2_data, branch_17_out1_data}), .valid_out_bus({branch_17_out2_valid, branch_17_out1_valid}), .ready_out_bus({branch_17_out2_ready, branch_17_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branch_18
		(.clk(branch_18_clk), .rst(branch_18_rst),
		.data_in_bus({{branch_18_in2_data}, branch_18_in1_data}), .valid_in_bus({branch_18_in2_valid, branch_18_in1_valid}), .ready_in_bus({branch_18_in2_ready, branch_18_in1_ready}), 
		.data_out_bus({branch_18_out2_data, branch_18_out1_data}), .valid_out_bus({branch_18_out2_valid, branch_18_out1_valid}), .ready_out_bus({branch_18_out2_ready, branch_18_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_33
		(.clk(fork_33_clk), .rst(fork_33_rst),
		.data_in_bus({fork_33_in1_data}), .valid_in_bus({fork_33_in1_valid}), .ready_in_bus({fork_33_in1_ready}), 
		.data_out_bus({fork_33_out4_data, fork_33_out3_data, fork_33_out2_data, fork_33_out1_data}), .valid_out_bus({fork_33_out4_valid, fork_33_out3_valid, fork_33_out2_valid, fork_33_out1_valid}), .ready_out_bus({fork_33_out4_ready, fork_33_out3_ready, fork_33_out2_ready, fork_33_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_35
		(.clk(phiC_35_clk), .rst(phiC_35_rst),
		.data_in_bus({phiC_35_in1_data}), .valid_in_bus({phiC_35_in1_valid}), .ready_in_bus({phiC_35_in1_ready}), 
		.data_out_bus({phiC_35_out1_data}), .valid_out_bus({phiC_35_out1_valid}), .ready_out_bus({phiC_35_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_48
		(.clk(forkC_48_clk), .rst(forkC_48_rst),
		.data_in_bus({forkC_48_in1_data}), .valid_in_bus({forkC_48_in1_valid}), .ready_in_bus({forkC_48_in1_ready}), 
		.data_out_bus({forkC_48_out5_data, forkC_48_out4_data, forkC_48_out3_data, forkC_48_out2_data, forkC_48_out1_data}), .valid_out_bus({forkC_48_out5_valid, forkC_48_out4_valid, forkC_48_out3_valid, forkC_48_out2_valid, forkC_48_out1_valid}), .ready_out_bus({forkC_48_out5_ready, forkC_48_out4_ready, forkC_48_out3_ready, forkC_48_out2_ready, forkC_48_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_50
		(.clk(branchC_50_clk), .rst(branchC_50_rst),
		.data_in_bus({{branchC_50_in2_data}, branchC_50_in1_data}), .valid_in_bus({branchC_50_in2_valid, branchC_50_in1_valid}), .ready_in_bus({branchC_50_in2_ready, branchC_50_in1_ready}), 
		.data_out_bus({branchC_50_out2_data, branchC_50_out1_data}), .valid_out_bus({branchC_50_out2_valid, branchC_50_out1_valid}), .ready_out_bus({branchC_50_out2_ready, branchC_50_out1_ready}));

	ret_op #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) ret_op_ret_0
		(.clk(ret_0_clk), .rst(ret_0_rst),
		.data_in_bus({ret_0_in1_data}), .valid_in_bus({ret_0_in1_valid}), .ready_in_bus({ret_0_in1_ready}), 
		.data_out_bus({ret_0_out1_data}), .valid_out_bus({ret_0_out1_valid}), .ready_out_bus({ret_0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n29
		(.clk(phi_n29_clk), .rst(phi_n29_rst),
		.data_in_bus({phi_n29_in1_data}), .valid_in_bus({phi_n29_in1_valid}), .ready_in_bus({phi_n29_in1_ready}), 
		.data_out_bus({phi_n29_out1_data}), .valid_out_bus({phi_n29_out1_valid}), .ready_out_bus({phi_n29_out1_ready}));

	end_node #(.INPUTS(1), .OUTPUTS(1), .MEMORY_INPUTS(3), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) end_node_end_0
		(.clk(end_0_clk), .rst(end_0_rst),
		.data_in_bus({end_0_in4_data}), .valid_in_bus({end_0_in4_valid}), .ready_in_bus({end_0_in4_ready}), .e_valid_bus({end_0_in3_valid, end_0_in2_valid, end_0_in1_valid}), .e_ready_bus({end_0_in3_ready, end_0_in2_ready, end_0_in1_ready}), 
		.data_out_bus({end_0_out1_data}), .valid_out_bus({end_0_out1_valid}), .ready_out_bus({end_0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_43
		(.clk(phiC_43_clk), .rst(phiC_43_rst),
		.data_in_bus({phiC_43_in1_data}), .valid_in_bus({phiC_43_in1_valid}), .ready_in_bus({phiC_43_in1_ready}), 
		.data_out_bus({phiC_43_out1_data}), .valid_out_bus({phiC_43_out1_valid}), .ready_out_bus({phiC_43_out1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_0
		(.clk(sink_0_clk), .rst(sink_0_rst),
		.data_in_bus({sink_0_in1_data}), .valid_in_bus({sink_0_in1_valid}), .ready_in_bus({sink_0_in1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_7
		(.clk(phi_7_clk), .rst(phi_7_rst),
		.data_in_bus({{31'b0, phi_7_in1_data}, phi_7_in3_data, phi_7_in2_data}), .valid_in_bus({phi_7_in1_valid, phi_7_in3_valid, phi_7_in2_valid}), .ready_in_bus({phi_7_in1_ready, phi_7_in3_ready, phi_7_in2_ready}), 
		.data_out_bus({phi_7_out1_data}), .valid_out_bus({phi_7_out1_valid}), .ready_out_bus({phi_7_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_3
		(.clk(cst_3_clk), .rst(cst_3_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_3_in1_valid}), .ready_in_bus({cst_3_in1_ready}), 
		.data_out_bus({cst_3_out1_data}), .valid_out_bus({cst_3_out1_valid}), .ready_out_bus({cst_3_out1_ready}));

	icmp_sgt_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(1)) icmp_sgt_op_icmp_8
		(.clk(icmp_8_clk), .rst(icmp_8_rst),
		.data_in_bus({icmp_8_in2_data, icmp_8_in1_data}), .valid_in_bus({icmp_8_in2_valid, icmp_8_in1_valid}), .ready_in_bus({icmp_8_in2_ready, icmp_8_in1_ready}), 
		.data_out_bus({icmp_8_out1_data}), .valid_out_bus({icmp_8_out1_valid}), .ready_out_bus({icmp_8_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n6
		(.clk(phi_n6_clk), .rst(phi_n6_rst),
		.data_in_bus({phi_n6_in2_data, phi_n6_in1_data}), .valid_in_bus({phi_n6_in2_valid, phi_n6_in1_valid}), .ready_in_bus({phi_n6_in2_ready, phi_n6_in1_ready}), 
		.data_out_bus({phi_n6_out1_data}), .valid_out_bus({phi_n6_out1_valid}), .ready_out_bus({phi_n6_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) merge_node_phi_n7
		(.clk(phi_n7_clk), .rst(phi_n7_rst),
		.data_in_bus({phi_n7_in2_data, phi_n7_in1_data}), .valid_in_bus({phi_n7_in2_valid, phi_n7_in1_valid}), .ready_in_bus({phi_n7_in2_ready, phi_n7_in1_ready}), 
		.data_out_bus({phi_n7_out1_data}), .valid_out_bus({phi_n7_out1_valid}), .ready_out_bus({phi_n7_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_1
		(.clk(fork_1_clk), .rst(fork_1_rst),
		.data_in_bus({fork_1_in1_data}), .valid_in_bus({fork_1_in1_valid}), .ready_in_bus({fork_1_in1_ready}), 
		.data_out_bus({fork_1_out2_data, fork_1_out1_data}), .valid_out_bus({fork_1_out2_valid, fork_1_out1_valid}), .ready_out_bus({fork_1_out2_ready, fork_1_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_5
		(.clk(branch_5_clk), .rst(branch_5_rst),
		.data_in_bus({{31'b0, branch_5_in2_data}, branch_5_in1_data}), .valid_in_bus({branch_5_in2_valid, branch_5_in1_valid}), .ready_in_bus({branch_5_in2_ready, branch_5_in1_ready}), 
		.data_out_bus({branch_5_out2_data, branch_5_out1_data}), .valid_out_bus({branch_5_out2_valid, branch_5_out1_valid}), .ready_out_bus({branch_5_out2_ready, branch_5_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_6
		(.clk(branch_6_clk), .rst(branch_6_rst),
		.data_in_bus({{31'b0, branch_6_in2_data}, branch_6_in1_data}), .valid_in_bus({branch_6_in2_valid, branch_6_in1_valid}), .ready_in_bus({branch_6_in2_ready, branch_6_in1_ready}), 
		.data_out_bus({branch_6_out2_data, branch_6_out1_data}), .valid_out_bus({branch_6_out2_valid, branch_6_out1_valid}), .ready_out_bus({branch_6_out2_ready, branch_6_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) branch_node_branch_7
		(.clk(branch_7_clk), .rst(branch_7_rst),
		.data_in_bus({{2'b0, branch_7_in2_data}, branch_7_in1_data}), .valid_in_bus({branch_7_in2_valid, branch_7_in1_valid}), .ready_in_bus({branch_7_in2_ready, branch_7_in1_ready}), 
		.data_out_bus({branch_7_out2_data, branch_7_out1_data}), .valid_out_bus({branch_7_out2_valid, branch_7_out1_valid}), .ready_out_bus({branch_7_out2_ready, branch_7_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_29
		(.clk(fork_29_clk), .rst(fork_29_rst),
		.data_in_bus({fork_29_in1_data}), .valid_in_bus({fork_29_in1_valid}), .ready_in_bus({fork_29_in1_ready}), 
		.data_out_bus({fork_29_out4_data, fork_29_out3_data, fork_29_out2_data, fork_29_out1_data}), .valid_out_bus({fork_29_out4_valid, fork_29_out3_valid, fork_29_out2_valid, fork_29_out1_valid}), .ready_out_bus({fork_29_out4_ready, fork_29_out3_ready, fork_29_out2_ready, fork_29_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_31
		(.clk(phiC_31_clk), .rst(phiC_31_rst),
		.data_in_bus({phiC_31_in2_data, phiC_31_in1_data}), .valid_in_bus({phiC_31_in2_valid, phiC_31_in1_valid}), .ready_in_bus({phiC_31_in2_ready, phiC_31_in1_ready}), 
		.data_out_bus({phiC_31_out2_data, phiC_31_out1_data}), .valid_out_bus({phiC_31_out2_valid, phiC_31_out1_valid}), .ready_out_bus({phiC_31_out2_ready, phiC_31_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_46
		(.clk(branchC_46_clk), .rst(branchC_46_rst),
		.data_in_bus({{branchC_46_in2_data}, branchC_46_in1_data}), .valid_in_bus({branchC_46_in2_valid, branchC_46_in1_valid}), .ready_in_bus({branchC_46_in2_ready, branchC_46_in1_ready}), 
		.data_out_bus({branchC_46_out2_data, branchC_46_out1_data}), .valid_out_bus({branchC_46_out2_valid, branchC_46_out1_valid}), .ready_out_bus({branchC_46_out2_ready, branchC_46_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_0
		(.clk(source_0_clk), .rst(source_0_rst),
		.data_out_bus({source_0_out1_data}), .valid_out_bus({source_0_out1_valid}), .ready_out_bus({source_0_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(3), .DATA_SIZE(32)) mc_load_op_load_17
		(.clk(load_17_clk), .rst(load_17_rst),
		.data_in_bus({load_17_in1_data}), .address_in_bus({load_17_in2_data}), .valid_in_bus({load_17_in2_valid, load_17_in1_valid}), .ready_in_bus({load_17_in2_ready, load_17_in1_ready}), 
		.data_out_bus({load_17_out1_data}), .address_out_bus({load_17_out2_data}), .valid_out_bus({load_17_out2_valid, load_17_out1_valid}), .ready_out_bus({load_17_out2_ready, load_17_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block5
		(.clk(brCst_block5_clk), .rst(brCst_block5_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block5_in1_valid}), .ready_in_bus({brCst_block5_in1_ready}), 
		.data_out_bus({brCst_block5_out1_data}), .valid_out_bus({brCst_block5_out1_valid}), .ready_out_bus({brCst_block5_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) merge_node_phi_n8
		(.clk(phi_n8_clk), .rst(phi_n8_rst),
		.data_in_bus({phi_n8_in1_data}), .valid_in_bus({phi_n8_in1_valid}), .ready_in_bus({phi_n8_in1_ready}), 
		.data_out_bus({phi_n8_out1_data}), .valid_out_bus({phi_n8_out1_valid}), .ready_out_bus({phi_n8_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n9
		(.clk(phi_n9_clk), .rst(phi_n9_rst),
		.data_in_bus({phi_n9_in1_data}), .valid_in_bus({phi_n9_in1_valid}), .ready_in_bus({phi_n9_in1_ready}), 
		.data_out_bus({phi_n9_out1_data}), .valid_out_bus({phi_n9_out1_valid}), .ready_out_bus({phi_n9_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) fork_node_fork_16
		(.clk(fork_16_clk), .rst(fork_16_rst),
		.data_in_bus({fork_16_in1_data}), .valid_in_bus({fork_16_in1_valid}), .ready_in_bus({fork_16_in1_ready}), 
		.data_out_bus({fork_16_out2_data, fork_16_out1_data}), .valid_out_bus({fork_16_out2_valid, fork_16_out1_valid}), .ready_out_bus({fork_16_out2_ready, fork_16_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_11
		(.clk(branch_11_clk), .rst(branch_11_rst),
		.data_in_bus({{31'b0, branch_11_in2_data}, branch_11_in1_data}), .valid_in_bus({branch_11_in2_valid, branch_11_in1_valid}), .ready_in_bus({branch_11_in2_ready, branch_11_in1_ready}), 
		.data_out_bus({branch_11_out2_data, branch_11_out1_data}), .valid_out_bus({branch_11_out2_valid, branch_11_out1_valid}), .ready_out_bus({branch_11_out2_ready, branch_11_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_12
		(.clk(branch_12_clk), .rst(branch_12_rst),
		.data_in_bus({{31'b0, branch_12_in2_data}, branch_12_in1_data}), .valid_in_bus({branch_12_in2_valid, branch_12_in1_valid}), .ready_in_bus({branch_12_in2_ready, branch_12_in1_ready}), 
		.data_out_bus({branch_12_out2_data, branch_12_out1_data}), .valid_out_bus({branch_12_out2_valid, branch_12_out1_valid}), .ready_out_bus({branch_12_out2_ready, branch_12_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) branch_node_branch_13
		(.clk(branch_13_clk), .rst(branch_13_rst),
		.data_in_bus({{2'b0, branch_13_in2_data}, branch_13_in1_data}), .valid_in_bus({branch_13_in2_valid, branch_13_in1_valid}), .ready_in_bus({branch_13_in2_ready, branch_13_in1_ready}), 
		.data_out_bus({branch_13_out2_data, branch_13_out1_data}), .valid_out_bus({branch_13_out2_valid, branch_13_out1_valid}), .ready_out_bus({branch_13_out2_ready, branch_13_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_31
		(.clk(fork_31_clk), .rst(fork_31_rst),
		.data_in_bus({fork_31_in1_data}), .valid_in_bus({fork_31_in1_valid}), .ready_in_bus({fork_31_in1_ready}), 
		.data_out_bus({fork_31_out4_data, fork_31_out3_data, fork_31_out2_data, fork_31_out1_data}), .valid_out_bus({fork_31_out4_valid, fork_31_out3_valid, fork_31_out2_valid, fork_31_out1_valid}), .ready_out_bus({fork_31_out4_ready, fork_31_out3_ready, fork_31_out2_ready, fork_31_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_33
		(.clk(phiC_33_clk), .rst(phiC_33_rst),
		.data_in_bus({phiC_33_in1_data}), .valid_in_bus({phiC_33_in1_valid}), .ready_in_bus({phiC_33_in1_ready}), 
		.data_out_bus({phiC_33_out1_data}), .valid_out_bus({phiC_33_out1_valid}), .ready_out_bus({phiC_33_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_46
		(.clk(forkC_46_clk), .rst(forkC_46_rst),
		.data_in_bus({forkC_46_in1_data}), .valid_in_bus({forkC_46_in1_valid}), .ready_in_bus({forkC_46_in1_ready}), 
		.data_out_bus({forkC_46_out2_data, forkC_46_out1_data}), .valid_out_bus({forkC_46_out2_valid, forkC_46_out1_valid}), .ready_out_bus({forkC_46_out2_ready, forkC_46_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_48
		(.clk(branchC_48_clk), .rst(branchC_48_rst),
		.data_in_bus({{branchC_48_in2_data}, branchC_48_in1_data}), .valid_in_bus({branchC_48_in2_valid, branchC_48_in1_valid}), .ready_in_bus({branchC_48_in2_ready, branchC_48_in1_ready}), 
		.data_out_bus({branchC_48_out2_data, branchC_48_out1_data}), .valid_out_bus({branchC_48_out2_valid, branchC_48_out1_valid}), .ready_out_bus({branchC_48_out2_ready, branchC_48_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_38
		(.clk(phi_38_clk), .rst(phi_38_rst),
		.data_in_bus({{31'b0, phi_38_in1_data}, phi_38_in3_data, phi_38_in2_data}), .valid_in_bus({phi_38_in1_valid, phi_38_in3_valid, phi_38_in2_valid}), .ready_in_bus({phi_38_in1_ready, phi_38_in3_ready, phi_38_in2_ready}), 
		.data_out_bus({phi_38_out1_data}), .valid_out_bus({phi_38_out1_valid}), .ready_out_bus({phi_38_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_9
		(.clk(cst_9_clk), .rst(cst_9_rst),
		.data_in_bus({1'd0}), .valid_in_bus({cst_9_in1_valid}), .ready_in_bus({cst_9_in1_ready}), 
		.data_out_bus({cst_9_out1_data}), .valid_out_bus({cst_9_out1_valid}), .ready_out_bus({cst_9_out1_ready}));

	icmp_sgt_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(1)) icmp_sgt_op_icmp_39
		(.clk(icmp_39_clk), .rst(icmp_39_rst),
		.data_in_bus({icmp_39_in2_data, icmp_39_in1_data}), .valid_in_bus({icmp_39_in2_valid, icmp_39_in1_valid}), .ready_in_bus({icmp_39_in2_ready, icmp_39_in1_ready}), 
		.data_out_bus({icmp_39_out1_data}), .valid_out_bus({icmp_39_out1_valid}), .ready_out_bus({icmp_39_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n10
		(.clk(phi_n10_clk), .rst(phi_n10_rst),
		.data_in_bus({phi_n10_in2_data, phi_n10_in1_data}), .valid_in_bus({phi_n10_in2_valid, phi_n10_in1_valid}), .ready_in_bus({phi_n10_in2_ready, phi_n10_in1_ready}), 
		.data_out_bus({phi_n10_out1_data}), .valid_out_bus({phi_n10_out1_valid}), .ready_out_bus({phi_n10_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n11
		(.clk(phi_n11_clk), .rst(phi_n11_rst),
		.data_in_bus({phi_n11_in2_data, phi_n11_in1_data}), .valid_in_bus({phi_n11_in2_valid, phi_n11_in1_valid}), .ready_in_bus({phi_n11_in2_ready, phi_n11_in1_ready}), 
		.data_out_bus({phi_n11_out1_data}), .valid_out_bus({phi_n11_out1_valid}), .ready_out_bus({phi_n11_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) merge_node_phi_n12
		(.clk(phi_n12_clk), .rst(phi_n12_rst),
		.data_in_bus({phi_n12_in2_data, phi_n12_in1_data}), .valid_in_bus({phi_n12_in2_valid, phi_n12_in1_valid}), .ready_in_bus({phi_n12_in2_ready, phi_n12_in1_ready}), 
		.data_out_bus({phi_n12_out1_data}), .valid_out_bus({phi_n12_out1_valid}), .ready_out_bus({phi_n12_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_5
		(.clk(fork_5_clk), .rst(fork_5_rst),
		.data_in_bus({fork_5_in1_data}), .valid_in_bus({fork_5_in1_valid}), .ready_in_bus({fork_5_in1_ready}), 
		.data_out_bus({fork_5_out2_data, fork_5_out1_data}), .valid_out_bus({fork_5_out2_valid, fork_5_out1_valid}), .ready_out_bus({fork_5_out2_ready, fork_5_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_23
		(.clk(branch_23_clk), .rst(branch_23_rst),
		.data_in_bus({{31'b0, branch_23_in2_data}, branch_23_in1_data}), .valid_in_bus({branch_23_in2_valid, branch_23_in1_valid}), .ready_in_bus({branch_23_in2_ready, branch_23_in1_ready}), 
		.data_out_bus({branch_23_out2_data, branch_23_out1_data}), .valid_out_bus({branch_23_out2_valid, branch_23_out1_valid}), .ready_out_bus({branch_23_out2_ready, branch_23_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_24
		(.clk(branch_24_clk), .rst(branch_24_rst),
		.data_in_bus({{31'b0, branch_24_in2_data}, branch_24_in1_data}), .valid_in_bus({branch_24_in2_valid, branch_24_in1_valid}), .ready_in_bus({branch_24_in2_ready, branch_24_in1_ready}), 
		.data_out_bus({branch_24_out2_data, branch_24_out1_data}), .valid_out_bus({branch_24_out2_valid, branch_24_out1_valid}), .ready_out_bus({branch_24_out2_ready, branch_24_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_25
		(.clk(branch_25_clk), .rst(branch_25_rst),
		.data_in_bus({{31'b0, branch_25_in2_data}, branch_25_in1_data}), .valid_in_bus({branch_25_in2_valid, branch_25_in1_valid}), .ready_in_bus({branch_25_in2_ready, branch_25_in1_ready}), 
		.data_out_bus({branch_25_out2_data, branch_25_out1_data}), .valid_out_bus({branch_25_out2_valid, branch_25_out1_valid}), .ready_out_bus({branch_25_out2_ready, branch_25_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) branch_node_branch_26
		(.clk(branch_26_clk), .rst(branch_26_rst),
		.data_in_bus({{9'b0, branch_26_in2_data}, branch_26_in1_data}), .valid_in_bus({branch_26_in2_valid, branch_26_in1_valid}), .ready_in_bus({branch_26_in2_ready, branch_26_in1_ready}), 
		.data_out_bus({branch_26_out2_data, branch_26_out1_data}), .valid_out_bus({branch_26_out2_valid, branch_26_out1_valid}), .ready_out_bus({branch_26_out2_ready, branch_26_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_35
		(.clk(fork_35_clk), .rst(fork_35_rst),
		.data_in_bus({fork_35_in1_data}), .valid_in_bus({fork_35_in1_valid}), .ready_in_bus({fork_35_in1_ready}), 
		.data_out_bus({fork_35_out5_data, fork_35_out4_data, fork_35_out3_data, fork_35_out2_data, fork_35_out1_data}), .valid_out_bus({fork_35_out5_valid, fork_35_out4_valid, fork_35_out3_valid, fork_35_out2_valid, fork_35_out1_valid}), .ready_out_bus({fork_35_out5_ready, fork_35_out4_ready, fork_35_out3_ready, fork_35_out2_ready, fork_35_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_37
		(.clk(phiC_37_clk), .rst(phiC_37_rst),
		.data_in_bus({phiC_37_in2_data, phiC_37_in1_data}), .valid_in_bus({phiC_37_in2_valid, phiC_37_in1_valid}), .ready_in_bus({phiC_37_in2_ready, phiC_37_in1_ready}), 
		.data_out_bus({phiC_37_out2_data, phiC_37_out1_data}), .valid_out_bus({phiC_37_out2_valid, phiC_37_out1_valid}), .ready_out_bus({phiC_37_out2_ready, phiC_37_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_52
		(.clk(branchC_52_clk), .rst(branchC_52_rst),
		.data_in_bus({{branchC_52_in2_data}, branchC_52_in1_data}), .valid_in_bus({branchC_52_in2_valid, branchC_52_in1_valid}), .ready_in_bus({branchC_52_in2_ready, branchC_52_in1_ready}), 
		.data_out_bus({branchC_52_out2_data, branchC_52_out1_data}), .valid_out_bus({branchC_52_out2_valid, branchC_52_out1_valid}), .ready_out_bus({branchC_52_out2_ready, branchC_52_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_3
		(.clk(source_3_clk), .rst(source_3_rst),
		.data_out_bus({source_3_out1_data}), .valid_out_bus({source_3_out1_valid}), .ready_out_bus({source_3_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(32), .DATA_SIZE(32)) mc_load_op_load_21
		(.clk(load_21_clk), .rst(load_21_rst),
		.data_in_bus({load_21_in1_data}), .address_in_bus({load_21_in2_data}), .valid_in_bus({load_21_in2_valid, load_21_in1_valid}), .ready_in_bus({load_21_in2_ready, load_21_in1_ready}), 
		.data_out_bus({load_21_out1_data}), .address_out_bus({load_21_out2_data}), .valid_out_bus({load_21_out2_valid, load_21_out1_valid}), .ready_out_bus({load_21_out2_ready, load_21_out1_ready}));

	icmp_eq_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(1)) icmp_eq_op_icmp_22
		(.clk(icmp_22_clk), .rst(icmp_22_rst),
		.data_in_bus({icmp_22_in2_data, icmp_22_in1_data}), .valid_in_bus({icmp_22_in2_valid, icmp_22_in1_valid}), .ready_in_bus({icmp_22_in2_ready, icmp_22_in1_ready}), 
		.data_out_bus({icmp_22_out1_data}), .valid_out_bus({icmp_22_out1_valid}), .ready_out_bus({icmp_22_out1_ready}));

	zext_op #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) zext_op_zext_23
		(.clk(zext_23_clk), .rst(zext_23_rst),
		.data_in_bus({zext_23_in1_data}), .valid_in_bus({zext_23_in1_valid}), .ready_in_bus({zext_23_in1_ready}), 
		.data_out_bus({zext_23_out1_data}), .valid_out_bus({zext_23_out1_valid}), .ready_out_bus({zext_23_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_24
		(.clk(add_24_clk), .rst(add_24_rst),
		.data_in_bus({add_24_in2_data, add_24_in1_data}), .valid_in_bus({add_24_in2_valid, add_24_in1_valid}), .ready_in_bus({add_24_in2_ready, add_24_in1_ready}), 
		.data_out_bus({add_24_out1_data}), .valid_out_bus({add_24_out1_valid}), .ready_out_bus({add_24_out1_ready}));

	mc_store_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(3), .DATA_SIZE(32)) mc_store_op_store_1
		(.clk(store_1_clk), .rst(store_1_rst),
		.data_in_bus({store_1_in1_data}), .address_in_bus({store_1_in2_data}), .valid_in_bus({store_1_in2_valid, store_1_in1_valid}), .ready_in_bus({store_1_in2_ready, store_1_in1_ready}), 
		.data_out_bus({store_1_out1_data}), .address_out_bus({store_1_out2_data}), .valid_out_bus({store_1_out2_valid, store_1_out1_valid}), .ready_out_bus({store_1_out2_ready, store_1_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_4
		(.clk(cst_4_clk), .rst(cst_4_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_4_in1_valid}), .ready_in_bus({cst_4_in1_ready}), 
		.data_out_bus({cst_4_out1_data}), .valid_out_bus({cst_4_out1_valid}), .ready_out_bus({cst_4_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) add_op_add_27
		(.clk(add_27_clk), .rst(add_27_rst),
		.data_in_bus({add_27_in2_data, add_27_in1_data}), .valid_in_bus({add_27_in2_valid, add_27_in1_valid}), .ready_in_bus({add_27_in2_ready, add_27_in1_ready}), 
		.data_out_bus({add_27_out1_data}), .valid_out_bus({add_27_out1_valid}), .ready_out_bus({add_27_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) const_node_cst_5
		(.clk(cst_5_clk), .rst(cst_5_rst),
		.data_in_bus({3'd4}), .valid_in_bus({cst_5_in1_valid}), .ready_in_bus({cst_5_in1_ready}), 
		.data_out_bus({cst_5_out1_data}), .valid_out_bus({cst_5_out1_valid}), .ready_out_bus({cst_5_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_28
		(.clk(icmp_28_clk), .rst(icmp_28_rst),
		.data_in_bus({icmp_28_in2_data, icmp_28_in1_data}), .valid_in_bus({icmp_28_in2_valid, icmp_28_in1_valid}), .ready_in_bus({icmp_28_in2_ready, icmp_28_in1_ready}), 
		.data_out_bus({icmp_28_out1_data}), .valid_out_bus({icmp_28_out1_valid}), .ready_out_bus({icmp_28_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n3
		(.clk(phi_n3_clk), .rst(phi_n3_rst),
		.data_in_bus({phi_n3_in2_data, phi_n3_in1_data}), .valid_in_bus({phi_n3_in2_valid, phi_n3_in1_valid}), .ready_in_bus({phi_n3_in2_ready, phi_n3_in1_ready}), 
		.data_out_bus({phi_n3_out1_data}), .valid_out_bus({phi_n3_out1_valid}), .ready_out_bus({phi_n3_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n4
		(.clk(phi_n4_clk), .rst(phi_n4_rst),
		.data_in_bus({phi_n4_in2_data, phi_n4_in1_data}), .valid_in_bus({phi_n4_in2_valid, phi_n4_in1_valid}), .ready_in_bus({phi_n4_in2_ready, phi_n4_in1_ready}), 
		.data_out_bus({phi_n4_out1_data}), .valid_out_bus({phi_n4_out1_valid}), .ready_out_bus({phi_n4_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) merge_node_phi_n5
		(.clk(phi_n5_clk), .rst(phi_n5_rst),
		.data_in_bus({phi_n5_in2_data, phi_n5_in1_data}), .valid_in_bus({phi_n5_in2_valid, phi_n5_in1_valid}), .ready_in_bus({phi_n5_in2_ready, phi_n5_in1_ready}), 
		.data_out_bus({phi_n5_out1_data}), .valid_out_bus({phi_n5_out1_valid}), .ready_out_bus({phi_n5_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_2
		(.clk(fork_2_clk), .rst(fork_2_rst),
		.data_in_bus({fork_2_in1_data}), .valid_in_bus({fork_2_in1_valid}), .ready_in_bus({fork_2_in1_ready}), 
		.data_out_bus({fork_2_out2_data, fork_2_out1_data}), .valid_out_bus({fork_2_out2_valid, fork_2_out1_valid}), .ready_out_bus({fork_2_out2_ready, fork_2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) fork_node_fork_3
		(.clk(fork_3_clk), .rst(fork_3_rst),
		.data_in_bus({fork_3_in1_data}), .valid_in_bus({fork_3_in1_valid}), .ready_in_bus({fork_3_in1_ready}), 
		.data_out_bus({fork_3_out2_data, fork_3_out1_data}), .valid_out_bus({fork_3_out2_valid, fork_3_out1_valid}), .ready_out_bus({fork_3_out2_ready, fork_3_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_12
		(.clk(fork_12_clk), .rst(fork_12_rst),
		.data_in_bus({fork_12_in1_data}), .valid_in_bus({fork_12_in1_valid}), .ready_in_bus({fork_12_in1_ready}), 
		.data_out_bus({fork_12_out2_data, fork_12_out1_data}), .valid_out_bus({fork_12_out2_valid, fork_12_out1_valid}), .ready_out_bus({fork_12_out2_ready, fork_12_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) fork_node_fork_13
		(.clk(fork_13_clk), .rst(fork_13_rst),
		.data_in_bus({fork_13_in1_data}), .valid_in_bus({fork_13_in1_valid}), .ready_in_bus({fork_13_in1_ready}), 
		.data_out_bus({fork_13_out2_data, fork_13_out1_data}), .valid_out_bus({fork_13_out2_valid, fork_13_out1_valid}), .ready_out_bus({fork_13_out2_ready, fork_13_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_14
		(.clk(branch_14_clk), .rst(branch_14_rst),
		.data_in_bus({{31'b0, branch_14_in2_data}, branch_14_in1_data}), .valid_in_bus({branch_14_in2_valid, branch_14_in1_valid}), .ready_in_bus({branch_14_in2_ready, branch_14_in1_ready}), 
		.data_out_bus({branch_14_out2_data, branch_14_out1_data}), .valid_out_bus({branch_14_out2_valid, branch_14_out1_valid}), .ready_out_bus({branch_14_out2_ready, branch_14_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) branch_node_branch_15
		(.clk(branch_15_clk), .rst(branch_15_rst),
		.data_in_bus({{2'b0, branch_15_in2_data}, branch_15_in1_data}), .valid_in_bus({branch_15_in2_valid, branch_15_in1_valid}), .ready_in_bus({branch_15_in2_ready, branch_15_in1_ready}), 
		.data_out_bus({branch_15_out2_data, branch_15_out1_data}), .valid_out_bus({branch_15_out2_valid, branch_15_out1_valid}), .ready_out_bus({branch_15_out2_ready, branch_15_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(3), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_32
		(.clk(fork_32_clk), .rst(fork_32_rst),
		.data_in_bus({fork_32_in1_data}), .valid_in_bus({fork_32_in1_valid}), .ready_in_bus({fork_32_in1_ready}), 
		.data_out_bus({fork_32_out3_data, fork_32_out2_data, fork_32_out1_data}), .valid_out_bus({fork_32_out3_valid, fork_32_out2_valid, fork_32_out1_valid}), .ready_out_bus({fork_32_out3_ready, fork_32_out2_ready, fork_32_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_17
		(.clk(cst_17_clk), .rst(cst_17_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_17_in1_valid}), .ready_in_bus({cst_17_in1_ready}), 
		.data_out_bus({cst_17_out1_data}), .valid_out_bus({cst_17_out1_valid}), .ready_out_bus({cst_17_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_34
		(.clk(phiC_34_clk), .rst(phiC_34_rst),
		.data_in_bus({phiC_34_in2_data, phiC_34_in1_data}), .valid_in_bus({phiC_34_in2_valid, phiC_34_in1_valid}), .ready_in_bus({phiC_34_in2_ready, phiC_34_in1_ready}), 
		.data_out_bus({phiC_34_out1_data}), .valid_out_bus({phiC_34_out1_valid}), .ready_out_bus({phiC_34_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_47
		(.clk(forkC_47_clk), .rst(forkC_47_rst),
		.data_in_bus({forkC_47_in1_data}), .valid_in_bus({forkC_47_in1_valid}), .ready_in_bus({forkC_47_in1_ready}), 
		.data_out_bus({forkC_47_out2_data, forkC_47_out1_data}), .valid_out_bus({forkC_47_out2_valid, forkC_47_out1_valid}), .ready_out_bus({forkC_47_out2_ready, forkC_47_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_49
		(.clk(branchC_49_clk), .rst(branchC_49_rst),
		.data_in_bus({{branchC_49_in2_data}, branchC_49_in1_data}), .valid_in_bus({branchC_49_in2_valid, branchC_49_in1_valid}), .ready_in_bus({branchC_49_in2_ready, branchC_49_in1_ready}), 
		.data_out_bus({branchC_49_out2_data, branchC_49_out1_data}), .valid_out_bus({branchC_49_out2_valid, branchC_49_out1_valid}), .ready_out_bus({branchC_49_out2_ready, branchC_49_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_1
		(.clk(source_1_clk), .rst(source_1_rst),
		.data_out_bus({source_1_out1_data}), .valid_out_bus({source_1_out1_valid}), .ready_out_bus({source_1_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(3))source_node_source_2
		(.clk(source_2_clk), .rst(source_2_rst),
		.data_out_bus({source_2_out1_data}), .valid_out_bus({source_2_out1_valid}), .ready_out_bus({source_2_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(32), .DATA_SIZE(32)) mc_load_op_load_12
		(.clk(load_12_clk), .rst(load_12_rst),
		.data_in_bus({load_12_in1_data}), .address_in_bus({load_12_in2_data}), .valid_in_bus({load_12_in2_valid, load_12_in1_valid}), .ready_in_bus({load_12_in2_ready, load_12_in1_ready}), 
		.data_out_bus({load_12_out1_data}), .address_out_bus({load_12_out2_data}), .valid_out_bus({load_12_out2_valid, load_12_out1_valid}), .ready_out_bus({load_12_out2_ready, load_12_out1_ready}));

	icmp_eq_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(1)) icmp_eq_op_icmp_13
		(.clk(icmp_13_clk), .rst(icmp_13_rst),
		.data_in_bus({icmp_13_in2_data, icmp_13_in1_data}), .valid_in_bus({icmp_13_in2_valid, icmp_13_in1_valid}), .ready_in_bus({icmp_13_in2_ready, icmp_13_in1_ready}), 
		.data_out_bus({icmp_13_out1_data}), .valid_out_bus({icmp_13_out1_valid}), .ready_out_bus({icmp_13_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n0
		(.clk(phi_n0_clk), .rst(phi_n0_rst),
		.data_in_bus({phi_n0_in1_data}), .valid_in_bus({phi_n0_in1_valid}), .ready_in_bus({phi_n0_in1_ready}), 
		.data_out_bus({phi_n0_out1_data}), .valid_out_bus({phi_n0_out1_valid}), .ready_out_bus({phi_n0_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n1
		(.clk(phi_n1_clk), .rst(phi_n1_rst),
		.data_in_bus({phi_n1_in1_data}), .valid_in_bus({phi_n1_in1_valid}), .ready_in_bus({phi_n1_in1_ready}), 
		.data_out_bus({phi_n1_out1_data}), .valid_out_bus({phi_n1_out1_valid}), .ready_out_bus({phi_n1_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) merge_node_phi_n2
		(.clk(phi_n2_clk), .rst(phi_n2_rst),
		.data_in_bus({phi_n2_in1_data}), .valid_in_bus({phi_n2_in1_valid}), .ready_in_bus({phi_n2_in1_ready}), 
		.data_out_bus({phi_n2_out1_data}), .valid_out_bus({phi_n2_out1_valid}), .ready_out_bus({phi_n2_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_9
		(.clk(fork_9_clk), .rst(fork_9_rst),
		.data_in_bus({fork_9_in1_data}), .valid_in_bus({fork_9_in1_valid}), .ready_in_bus({fork_9_in1_ready}), 
		.data_out_bus({fork_9_out2_data, fork_9_out1_data}), .valid_out_bus({fork_9_out2_valid, fork_9_out1_valid}), .ready_out_bus({fork_9_out2_ready, fork_9_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_10
		(.clk(fork_10_clk), .rst(fork_10_rst),
		.data_in_bus({fork_10_in1_data}), .valid_in_bus({fork_10_in1_valid}), .ready_in_bus({fork_10_in1_ready}), 
		.data_out_bus({fork_10_out2_data, fork_10_out1_data}), .valid_out_bus({fork_10_out2_valid, fork_10_out1_valid}), .ready_out_bus({fork_10_out2_ready, fork_10_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_8
		(.clk(branch_8_clk), .rst(branch_8_rst),
		.data_in_bus({{31'b0, branch_8_in2_data}, branch_8_in1_data}), .valid_in_bus({branch_8_in2_valid, branch_8_in1_valid}), .ready_in_bus({branch_8_in2_ready, branch_8_in1_ready}), 
		.data_out_bus({branch_8_out2_data, branch_8_out1_data}), .valid_out_bus({branch_8_out2_valid, branch_8_out1_valid}), .ready_out_bus({branch_8_out2_ready, branch_8_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_9
		(.clk(branch_9_clk), .rst(branch_9_rst),
		.data_in_bus({{31'b0, branch_9_in2_data}, branch_9_in1_data}), .valid_in_bus({branch_9_in2_valid, branch_9_in1_valid}), .ready_in_bus({branch_9_in2_ready, branch_9_in1_ready}), 
		.data_out_bus({branch_9_out2_data, branch_9_out1_data}), .valid_out_bus({branch_9_out2_valid, branch_9_out1_valid}), .ready_out_bus({branch_9_out2_ready, branch_9_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(3), .DATA_OUT_SIZE(3)) branch_node_branch_10
		(.clk(branch_10_clk), .rst(branch_10_rst),
		.data_in_bus({{2'b0, branch_10_in2_data}, branch_10_in1_data}), .valid_in_bus({branch_10_in2_valid, branch_10_in1_valid}), .ready_in_bus({branch_10_in2_ready, branch_10_in1_ready}), 
		.data_out_bus({branch_10_out2_data, branch_10_out1_data}), .valid_out_bus({branch_10_out2_valid, branch_10_out1_valid}), .ready_out_bus({branch_10_out2_ready, branch_10_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_30
		(.clk(fork_30_clk), .rst(fork_30_rst),
		.data_in_bus({fork_30_in1_data}), .valid_in_bus({fork_30_in1_valid}), .ready_in_bus({fork_30_in1_ready}), 
		.data_out_bus({fork_30_out4_data, fork_30_out3_data, fork_30_out2_data, fork_30_out1_data}), .valid_out_bus({fork_30_out4_valid, fork_30_out3_valid, fork_30_out2_valid, fork_30_out1_valid}), .ready_out_bus({fork_30_out4_ready, fork_30_out3_ready, fork_30_out2_ready, fork_30_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_32
		(.clk(phiC_32_clk), .rst(phiC_32_rst),
		.data_in_bus({phiC_32_in1_data}), .valid_in_bus({phiC_32_in1_valid}), .ready_in_bus({phiC_32_in1_ready}), 
		.data_out_bus({phiC_32_out1_data}), .valid_out_bus({phiC_32_out1_valid}), .ready_out_bus({phiC_32_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_47
		(.clk(branchC_47_clk), .rst(branchC_47_rst),
		.data_in_bus({{branchC_47_in2_data}, branchC_47_in1_data}), .valid_in_bus({branchC_47_in2_valid, branchC_47_in1_valid}), .ready_in_bus({branchC_47_in2_ready, branchC_47_in1_ready}), 
		.data_out_bus({branchC_47_out2_data, branchC_47_out1_data}), .valid_out_bus({branchC_47_out2_valid, branchC_47_out1_valid}), .ready_out_bus({branchC_47_out2_ready, branchC_47_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_64
		(.clk(phi_64_clk), .rst(phi_64_rst),
		.data_in_bus({{31'b0, phi_64_in1_data}, phi_64_in3_data, phi_64_in2_data}), .valid_in_bus({phi_64_in1_valid, phi_64_in3_valid, phi_64_in2_valid}), .ready_in_bus({phi_64_in1_ready, phi_64_in3_ready, phi_64_in2_ready}), 
		.data_out_bus({phi_64_out1_data}), .valid_out_bus({phi_64_out1_valid}), .ready_out_bus({phi_64_out1_ready}));

	mux_node #(.INPUTS(3), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32), .COND_SIZE(1)) mux_node_phi_65
		(.clk(phi_65_clk), .rst(phi_65_rst),
		.data_in_bus({{31'b0, phi_65_in1_data}, phi_65_in3_data, phi_65_in2_data}), .valid_in_bus({phi_65_in1_valid, phi_65_in3_valid, phi_65_in2_valid}), .ready_in_bus({phi_65_in1_ready, phi_65_in3_ready, phi_65_in2_ready}), 
		.data_out_bus({phi_65_out1_data}), .valid_out_bus({phi_65_out1_valid}), .ready_out_bus({phi_65_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_13
		(.clk(cst_13_clk), .rst(cst_13_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_13_in1_valid}), .ready_in_bus({cst_13_in1_ready}), 
		.data_out_bus({cst_13_out1_data}), .valid_out_bus({cst_13_out1_valid}), .ready_out_bus({cst_13_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) add_op_add_66
		(.clk(add_66_clk), .rst(add_66_rst),
		.data_in_bus({add_66_in2_data, add_66_in1_data}), .valid_in_bus({add_66_in2_valid, add_66_in1_valid}), .ready_in_bus({add_66_in2_ready, add_66_in1_ready}), 
		.data_out_bus({add_66_out1_data}), .valid_out_bus({add_66_out1_valid}), .ready_out_bus({add_66_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) const_node_cst_14
		(.clk(cst_14_clk), .rst(cst_14_rst),
		.data_in_bus({10'd1000}), .valid_in_bus({cst_14_in1_valid}), .ready_in_bus({cst_14_in1_ready}), 
		.data_out_bus({cst_14_out1_data}), .valid_out_bus({cst_14_out1_valid}), .ready_out_bus({cst_14_out1_ready}));

	icmp_ult_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(1)) icmp_ult_op_icmp_67
		(.clk(icmp_67_clk), .rst(icmp_67_rst),
		.data_in_bus({icmp_67_in2_data, icmp_67_in1_data}), .valid_in_bus({icmp_67_in2_valid, icmp_67_in1_valid}), .ready_in_bus({icmp_67_in2_ready, icmp_67_in1_ready}), 
		.data_out_bus({icmp_67_out1_data}), .valid_out_bus({icmp_67_out1_valid}), .ready_out_bus({icmp_67_out1_ready}));

	merge_node #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) merge_node_phi_n16
		(.clk(phi_n16_clk), .rst(phi_n16_rst),
		.data_in_bus({phi_n16_in2_data, phi_n16_in1_data}), .valid_in_bus({phi_n16_in2_valid, phi_n16_in1_valid}), .ready_in_bus({phi_n16_in2_ready, phi_n16_in1_ready}), 
		.data_out_bus({phi_n16_out1_data}), .valid_out_bus({phi_n16_out1_valid}), .ready_out_bus({phi_n16_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) fork_node_fork_8
		(.clk(fork_8_clk), .rst(fork_8_rst),
		.data_in_bus({fork_8_in1_data}), .valid_in_bus({fork_8_in1_valid}), .ready_in_bus({fork_8_in1_ready}), 
		.data_out_bus({fork_8_out2_data, fork_8_out1_data}), .valid_out_bus({fork_8_out2_valid, fork_8_out1_valid}), .ready_out_bus({fork_8_out2_ready, fork_8_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_41
		(.clk(branch_41_clk), .rst(branch_41_rst),
		.data_in_bus({{31'b0, branch_41_in2_data}, branch_41_in1_data}), .valid_in_bus({branch_41_in2_valid, branch_41_in1_valid}), .ready_in_bus({branch_41_in2_ready, branch_41_in1_ready}), 
		.data_out_bus({branch_41_out2_data, branch_41_out1_data}), .valid_out_bus({branch_41_out2_valid, branch_41_out1_valid}), .ready_out_bus({branch_41_out2_ready, branch_41_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_42
		(.clk(branch_42_clk), .rst(branch_42_rst),
		.data_in_bus({{31'b0, branch_42_in2_data}, branch_42_in1_data}), .valid_in_bus({branch_42_in2_valid, branch_42_in1_valid}), .ready_in_bus({branch_42_in2_ready, branch_42_in1_ready}), 
		.data_out_bus({branch_42_out2_data, branch_42_out1_data}), .valid_out_bus({branch_42_out2_valid, branch_42_out1_valid}), .ready_out_bus({branch_42_out2_ready, branch_42_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) branch_node_branch_43
		(.clk(branch_43_clk), .rst(branch_43_rst),
		.data_in_bus({{9'b0, branch_43_in2_data}, branch_43_in1_data}), .valid_in_bus({branch_43_in2_valid, branch_43_in1_valid}), .ready_in_bus({branch_43_in2_ready, branch_43_in1_ready}), 
		.data_out_bus({branch_43_out2_data, branch_43_out1_data}), .valid_out_bus({branch_43_out2_valid, branch_43_out1_valid}), .ready_out_bus({branch_43_out2_ready, branch_43_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_40
		(.clk(fork_40_clk), .rst(fork_40_rst),
		.data_in_bus({fork_40_in1_data}), .valid_in_bus({fork_40_in1_valid}), .ready_in_bus({fork_40_in1_ready}), 
		.data_out_bus({fork_40_out4_data, fork_40_out3_data, fork_40_out2_data, fork_40_out1_data}), .valid_out_bus({fork_40_out4_valid, fork_40_out3_valid, fork_40_out2_valid, fork_40_out1_valid}), .ready_out_bus({fork_40_out4_ready, fork_40_out3_ready, fork_40_out2_ready, fork_40_out1_ready}));

	cntrlMerge_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) cntrlMerge_node_phiC_42
		(.clk(phiC_42_clk), .rst(phiC_42_rst),
		.data_in_bus({phiC_42_in2_data, phiC_42_in1_data}), .valid_in_bus({phiC_42_in2_valid, phiC_42_in1_valid}), .ready_in_bus({phiC_42_in2_ready, phiC_42_in1_ready}), 
		.data_out_bus({phiC_42_out2_data, phiC_42_out1_data}), .valid_out_bus({phiC_42_out2_valid, phiC_42_out1_valid}), .ready_out_bus({phiC_42_out2_ready, phiC_42_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_57
		(.clk(branchC_57_clk), .rst(branchC_57_rst),
		.data_in_bus({{branchC_57_in2_data}, branchC_57_in1_data}), .valid_in_bus({branchC_57_in2_valid, branchC_57_in1_valid}), .ready_in_bus({branchC_57_in2_ready, branchC_57_in1_ready}), 
		.data_out_bus({branchC_57_out2_data, branchC_57_out1_data}), .valid_out_bus({branchC_57_out2_valid, branchC_57_out1_valid}), .ready_out_bus({branchC_57_out2_ready, branchC_57_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_7
		(.clk(source_7_clk), .rst(source_7_rst),
		.data_out_bus({source_7_out1_data}), .valid_out_bus({source_7_out1_valid}), .ready_out_bus({source_7_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(10))source_node_source_8
		(.clk(source_8_clk), .rst(source_8_rst),
		.data_out_bus({source_8_out1_data}), .valid_out_bus({source_8_out1_valid}), .ready_out_bus({source_8_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_61
		(.clk(fork_61_clk), .rst(fork_61_rst),
		.data_in_bus({fork_61_in1_data}), .valid_in_bus({fork_61_in1_valid}), .ready_in_bus({fork_61_in1_ready}), 
		.data_out_bus({fork_61_out2_data, fork_61_out1_data}), .valid_out_bus({fork_61_out2_valid, fork_61_out1_valid}), .ready_out_bus({fork_61_out2_ready, fork_61_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_cst_11
		(.clk(cst_11_clk), .rst(cst_11_rst),
		.data_in_bus({1'd1}), .valid_in_bus({cst_11_in1_valid}), .ready_in_bus({cst_11_in1_ready}), 
		.data_out_bus({cst_11_out1_data}), .valid_out_bus({cst_11_out1_valid}), .ready_out_bus({cst_11_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_58
		(.clk(add_58_clk), .rst(add_58_rst),
		.data_in_bus({add_58_in2_data, add_58_in1_data}), .valid_in_bus({add_58_in2_valid, add_58_in1_valid}), .ready_in_bus({add_58_in2_ready, add_58_in1_ready}), 
		.data_out_bus({add_58_out1_data}), .valid_out_bus({add_58_out1_valid}), .ready_out_bus({add_58_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) const_node_cst_12
		(.clk(cst_12_clk), .rst(cst_12_rst),
		.data_in_bus({32'd4294967295}), .valid_in_bus({cst_12_in1_valid}), .ready_in_bus({cst_12_in1_ready}), 
		.data_out_bus({cst_12_out1_data}), .valid_out_bus({cst_12_out1_valid}), .ready_out_bus({cst_12_out1_ready}));

	add_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) add_op_add_59
		(.clk(add_59_clk), .rst(add_59_rst),
		.data_in_bus({add_59_in2_data, add_59_in1_data}), .valid_in_bus({add_59_in2_valid, add_59_in1_valid}), .ready_in_bus({add_59_in2_ready, add_59_in1_ready}), 
		.data_out_bus({add_59_out1_data}), .valid_out_bus({add_59_out1_valid}), .ready_out_bus({add_59_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(32), .DATA_SIZE(32)) mc_load_op_load_62
		(.clk(load_62_clk), .rst(load_62_rst),
		.data_in_bus({load_62_in1_data}), .address_in_bus({load_62_in2_data}), .valid_in_bus({load_62_in2_valid, load_62_in1_valid}), .ready_in_bus({load_62_in2_ready, load_62_in1_ready}), 
		.data_out_bus({load_62_out1_data}), .address_out_bus({load_62_out2_data}), .valid_out_bus({load_62_out2_valid, load_62_out1_valid}), .ready_out_bus({load_62_out2_ready, load_62_out1_ready}));

	const_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) const_node_brCst_block13
		(.clk(brCst_block13_clk), .rst(brCst_block13_rst),
		.data_in_bus({1'd1}), .valid_in_bus({brCst_block13_in1_valid}), .ready_in_bus({brCst_block13_in1_ready}), 
		.data_out_bus({brCst_block13_out1_data}), .valid_out_bus({brCst_block13_out1_valid}), .ready_out_bus({brCst_block13_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n13
		(.clk(phi_n13_clk), .rst(phi_n13_rst),
		.data_in_bus({phi_n13_in1_data}), .valid_in_bus({phi_n13_in1_valid}), .ready_in_bus({phi_n13_in1_ready}), 
		.data_out_bus({phi_n13_out1_data}), .valid_out_bus({phi_n13_out1_valid}), .ready_out_bus({phi_n13_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n14
		(.clk(phi_n14_clk), .rst(phi_n14_rst),
		.data_in_bus({phi_n14_in1_data}), .valid_in_bus({phi_n14_in1_valid}), .ready_in_bus({phi_n14_in1_ready}), 
		.data_out_bus({phi_n14_out1_data}), .valid_out_bus({phi_n14_out1_valid}), .ready_out_bus({phi_n14_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) merge_node_phi_n15
		(.clk(phi_n15_clk), .rst(phi_n15_rst),
		.data_in_bus({phi_n15_in1_data}), .valid_in_bus({phi_n15_in1_valid}), .ready_in_bus({phi_n15_in1_ready}), 
		.data_out_bus({phi_n15_out1_data}), .valid_out_bus({phi_n15_out1_valid}), .ready_out_bus({phi_n15_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_38
		(.clk(branch_38_clk), .rst(branch_38_rst),
		.data_in_bus({{31'b0, branch_38_in2_data}, branch_38_in1_data}), .valid_in_bus({branch_38_in2_valid, branch_38_in1_valid}), .ready_in_bus({branch_38_in2_ready, branch_38_in1_ready}), 
		.data_out_bus({branch_38_out2_data, branch_38_out1_data}), .valid_out_bus({branch_38_out2_valid, branch_38_out1_valid}), .ready_out_bus({branch_38_out2_ready, branch_38_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_39
		(.clk(branch_39_clk), .rst(branch_39_rst),
		.data_in_bus({{31'b0, branch_39_in2_data}, branch_39_in1_data}), .valid_in_bus({branch_39_in2_valid, branch_39_in1_valid}), .ready_in_bus({branch_39_in2_ready, branch_39_in1_ready}), 
		.data_out_bus({branch_39_out2_data, branch_39_out1_data}), .valid_out_bus({branch_39_out2_valid, branch_39_out1_valid}), .ready_out_bus({branch_39_out2_ready, branch_39_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) branch_node_branch_40
		(.clk(branch_40_clk), .rst(branch_40_rst),
		.data_in_bus({{9'b0, branch_40_in2_data}, branch_40_in1_data}), .valid_in_bus({branch_40_in2_valid, branch_40_in1_valid}), .ready_in_bus({branch_40_in2_ready, branch_40_in1_ready}), 
		.data_out_bus({branch_40_out2_data, branch_40_out1_data}), .valid_out_bus({branch_40_out2_valid, branch_40_out1_valid}), .ready_out_bus({branch_40_out2_ready, branch_40_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(4), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_39
		(.clk(fork_39_clk), .rst(fork_39_rst),
		.data_in_bus({fork_39_in1_data}), .valid_in_bus({fork_39_in1_valid}), .ready_in_bus({fork_39_in1_ready}), 
		.data_out_bus({fork_39_out4_data, fork_39_out3_data, fork_39_out2_data, fork_39_out1_data}), .valid_out_bus({fork_39_out4_valid, fork_39_out3_valid, fork_39_out2_valid, fork_39_out1_valid}), .ready_out_bus({fork_39_out4_ready, fork_39_out3_ready, fork_39_out2_ready, fork_39_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_41
		(.clk(phiC_41_clk), .rst(phiC_41_rst),
		.data_in_bus({phiC_41_in1_data}), .valid_in_bus({phiC_41_in1_valid}), .ready_in_bus({phiC_41_in1_ready}), 
		.data_out_bus({phiC_41_out1_data}), .valid_out_bus({phiC_41_out1_valid}), .ready_out_bus({phiC_41_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_forkC_54
		(.clk(forkC_54_clk), .rst(forkC_54_rst),
		.data_in_bus({forkC_54_in1_data}), .valid_in_bus({forkC_54_in1_valid}), .ready_in_bus({forkC_54_in1_ready}), 
		.data_out_bus({forkC_54_out2_data, forkC_54_out1_data}), .valid_out_bus({forkC_54_out2_valid, forkC_54_out1_valid}), .ready_out_bus({forkC_54_out2_ready, forkC_54_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_56
		(.clk(branchC_56_clk), .rst(branchC_56_rst),
		.data_in_bus({{branchC_56_in2_data}, branchC_56_in1_data}), .valid_in_bus({branchC_56_in2_valid, branchC_56_in1_valid}), .ready_in_bus({branchC_56_in2_ready, branchC_56_in1_ready}), 
		.data_out_bus({branchC_56_out2_data, branchC_56_out1_data}), .valid_out_bus({branchC_56_out2_valid, branchC_56_out1_valid}), .ready_out_bus({branchC_56_out2_ready, branchC_56_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(1))source_node_source_5
		(.clk(source_5_clk), .rst(source_5_rst),
		.data_out_bus({source_5_out1_data}), .valid_out_bus({source_5_out1_valid}), .ready_out_bus({source_5_out1_ready}));

	source_node #(.INPUTS(0), .OUTPUTS(1), .DATA_OUT_SIZE(32))source_node_source_6
		(.clk(source_6_clk), .rst(source_6_rst),
		.data_out_bus({source_6_out1_data}), .valid_out_bus({source_6_out1_valid}), .ready_out_bus({source_6_out1_ready}));

	mc_load_op #(.INPUTS(2), .OUTPUTS(2), .ADDRESS_SIZE(32), .DATA_SIZE(32)) mc_load_op_load_43
		(.clk(load_43_clk), .rst(load_43_rst),
		.data_in_bus({load_43_in1_data}), .address_in_bus({load_43_in2_data}), .valid_in_bus({load_43_in2_valid, load_43_in1_valid}), .ready_in_bus({load_43_in2_ready, load_43_in1_ready}), 
		.data_out_bus({load_43_out1_data}), .address_out_bus({load_43_out2_data}), .valid_out_bus({load_43_out2_valid, load_43_out1_valid}), .ready_out_bus({load_43_out2_ready, load_43_out1_ready}));

	icmp_eq_op #(.INPUTS(2), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(1)) icmp_eq_op_icmp_44
		(.clk(icmp_44_clk), .rst(icmp_44_rst),
		.data_in_bus({icmp_44_in2_data, icmp_44_in1_data}), .valid_in_bus({icmp_44_in2_valid, icmp_44_in1_valid}), .ready_in_bus({icmp_44_in2_ready, icmp_44_in1_ready}), 
		.data_out_bus({icmp_44_out1_data}), .valid_out_bus({icmp_44_out1_valid}), .ready_out_bus({icmp_44_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n21
		(.clk(phi_n21_clk), .rst(phi_n21_rst),
		.data_in_bus({phi_n21_in1_data}), .valid_in_bus({phi_n21_in1_valid}), .ready_in_bus({phi_n21_in1_ready}), 
		.data_out_bus({phi_n21_out1_data}), .valid_out_bus({phi_n21_out1_valid}), .ready_out_bus({phi_n21_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n22
		(.clk(phi_n22_clk), .rst(phi_n22_rst),
		.data_in_bus({phi_n22_in1_data}), .valid_in_bus({phi_n22_in1_valid}), .ready_in_bus({phi_n22_in1_ready}), 
		.data_out_bus({phi_n22_out1_data}), .valid_out_bus({phi_n22_out1_valid}), .ready_out_bus({phi_n22_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) merge_node_phi_n23
		(.clk(phi_n23_clk), .rst(phi_n23_rst),
		.data_in_bus({phi_n23_in1_data}), .valid_in_bus({phi_n23_in1_valid}), .ready_in_bus({phi_n23_in1_ready}), 
		.data_out_bus({phi_n23_out1_data}), .valid_out_bus({phi_n23_out1_valid}), .ready_out_bus({phi_n23_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) merge_node_phi_n24
		(.clk(phi_n24_clk), .rst(phi_n24_rst),
		.data_in_bus({phi_n24_in1_data}), .valid_in_bus({phi_n24_in1_valid}), .ready_in_bus({phi_n24_in1_ready}), 
		.data_out_bus({phi_n24_out1_data}), .valid_out_bus({phi_n24_out1_valid}), .ready_out_bus({phi_n24_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_20
		(.clk(fork_20_clk), .rst(fork_20_rst),
		.data_in_bus({fork_20_in1_data}), .valid_in_bus({fork_20_in1_valid}), .ready_in_bus({fork_20_in1_ready}), 
		.data_out_bus({fork_20_out2_data, fork_20_out1_data}), .valid_out_bus({fork_20_out2_valid, fork_20_out1_valid}), .ready_out_bus({fork_20_out2_ready, fork_20_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) fork_node_fork_21
		(.clk(fork_21_clk), .rst(fork_21_rst),
		.data_in_bus({fork_21_in1_data}), .valid_in_bus({fork_21_in1_valid}), .ready_in_bus({fork_21_in1_ready}), 
		.data_out_bus({fork_21_out2_data, fork_21_out1_data}), .valid_out_bus({fork_21_out2_valid, fork_21_out1_valid}), .ready_out_bus({fork_21_out2_ready, fork_21_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_27
		(.clk(branch_27_clk), .rst(branch_27_rst),
		.data_in_bus({{31'b0, branch_27_in2_data}, branch_27_in1_data}), .valid_in_bus({branch_27_in2_valid, branch_27_in1_valid}), .ready_in_bus({branch_27_in2_ready, branch_27_in1_ready}), 
		.data_out_bus({branch_27_out2_data, branch_27_out1_data}), .valid_out_bus({branch_27_out2_valid, branch_27_out1_valid}), .ready_out_bus({branch_27_out2_ready, branch_27_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_28
		(.clk(branch_28_clk), .rst(branch_28_rst),
		.data_in_bus({{31'b0, branch_28_in2_data}, branch_28_in1_data}), .valid_in_bus({branch_28_in2_valid, branch_28_in1_valid}), .ready_in_bus({branch_28_in2_ready, branch_28_in1_ready}), 
		.data_out_bus({branch_28_out2_data, branch_28_out1_data}), .valid_out_bus({branch_28_out2_valid, branch_28_out1_valid}), .ready_out_bus({branch_28_out2_ready, branch_28_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) branch_node_branch_29
		(.clk(branch_29_clk), .rst(branch_29_rst),
		.data_in_bus({{31'b0, branch_29_in2_data}, branch_29_in1_data}), .valid_in_bus({branch_29_in2_valid, branch_29_in1_valid}), .ready_in_bus({branch_29_in2_ready, branch_29_in1_ready}), 
		.data_out_bus({branch_29_out2_data, branch_29_out1_data}), .valid_out_bus({branch_29_out2_valid, branch_29_out1_valid}), .ready_out_bus({branch_29_out2_ready, branch_29_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(10), .DATA_OUT_SIZE(10)) branch_node_branch_30
		(.clk(branch_30_clk), .rst(branch_30_rst),
		.data_in_bus({{9'b0, branch_30_in2_data}, branch_30_in1_data}), .valid_in_bus({branch_30_in2_valid, branch_30_in1_valid}), .ready_in_bus({branch_30_in2_ready, branch_30_in1_ready}), 
		.data_out_bus({branch_30_out2_data, branch_30_out1_data}), .valid_out_bus({branch_30_out2_valid, branch_30_out1_valid}), .ready_out_bus({branch_30_out2_ready, branch_30_out1_ready}));

	fork_node #(.INPUTS(1), .OUTPUTS(5), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) fork_node_fork_36
		(.clk(fork_36_clk), .rst(fork_36_rst),
		.data_in_bus({fork_36_in1_data}), .valid_in_bus({fork_36_in1_valid}), .ready_in_bus({fork_36_in1_ready}), 
		.data_out_bus({fork_36_out5_data, fork_36_out4_data, fork_36_out3_data, fork_36_out2_data, fork_36_out1_data}), .valid_out_bus({fork_36_out5_valid, fork_36_out4_valid, fork_36_out3_valid, fork_36_out2_valid, fork_36_out1_valid}), .ready_out_bus({fork_36_out5_ready, fork_36_out4_ready, fork_36_out3_ready, fork_36_out2_ready, fork_36_out1_ready}));

	merge_node #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) merge_node_phiC_38
		(.clk(phiC_38_clk), .rst(phiC_38_rst),
		.data_in_bus({phiC_38_in1_data}), .valid_in_bus({phiC_38_in1_valid}), .ready_in_bus({phiC_38_in1_ready}), 
		.data_out_bus({phiC_38_out1_data}), .valid_out_bus({phiC_38_out1_valid}), .ready_out_bus({phiC_38_out1_ready}));

	branch_node #(.INPUTS(2), .OUTPUTS(2), .DATA_IN_SIZE(1), .DATA_OUT_SIZE(1)) branch_node_branchC_53
		(.clk(branchC_53_clk), .rst(branchC_53_rst),
		.data_in_bus({{branchC_53_in2_data}, branchC_53_in1_data}), .valid_in_bus({branchC_53_in2_valid, branchC_53_in1_valid}), .ready_in_bus({branchC_53_in2_ready, branchC_53_in1_ready}), 
		.data_out_bus({branchC_53_out2_data, branchC_53_out1_data}), .valid_out_bus({branchC_53_out2_valid, branchC_53_out1_valid}), .ready_out_bus({branchC_53_out2_ready, branchC_53_out1_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(32), .BB_COUNT(2), .LOAD_COUNT(3), .STORE_COUNT(2))MemCont_MC_kmpNext
		(.clk(MC_kmpNext_clk), .rst(MC_kmpNext_rst),
		.io_storeDataOut(kmpNext_dout0), .io_storeAddrOut(kmpNext_address0), .io_storeEnable(kmpNext_we0),
		.io_loadDataIn(kmpNext_din1), .io_loadAddrOut(kmpNext_address1), .io_loadEnable(kmpNext_ce1),
		.io_bbpValids({MC_kmpNext_in2_valid, MC_kmpNext_in1_valid}), .io_bb_stCountArray({MC_kmpNext_in2_data, MC_kmpNext_in1_data}), .io_bbReadyToPrevs({MC_kmpNext_in2_ready, MC_kmpNext_in1_ready}), .io_rdPortsPrev_ready({MC_kmpNext_in9_ready, MC_kmpNext_in8_ready, MC_kmpNext_in5_ready}), .io_rdPortsPrev_valid({MC_kmpNext_in9_valid, MC_kmpNext_in8_valid, MC_kmpNext_in5_valid}), .io_rdPortsPrev_bits({MC_kmpNext_in9_data, MC_kmpNext_in8_data, MC_kmpNext_in5_data}), 	
	.io_wrAddrPorts_ready({MC_kmpNext_in6_ready, MC_kmpNext_in3_ready}), .io_wrAddrPorts_valid({MC_kmpNext_in6_valid, MC_kmpNext_in3_valid}), .io_wrAddrPorts_bits({MC_kmpNext_in6_data, MC_kmpNext_in3_data}), 	
	.io_wrDataPorts_ready({MC_kmpNext_in7_ready, MC_kmpNext_in4_ready}), .io_wrDataPorts_valid({MC_kmpNext_in7_valid, MC_kmpNext_in4_valid}), .io_wrDataPorts_bits({MC_kmpNext_in7_data, MC_kmpNext_in4_data}), 	
	.io_rdPortsNext_ready({MC_kmpNext_out3_ready, MC_kmpNext_out2_ready, MC_kmpNext_out1_ready}), .io_rdPortsNext_valid({MC_kmpNext_out3_valid, MC_kmpNext_out2_valid, MC_kmpNext_out1_valid}), .io_rdPortsNext_bits({MC_kmpNext_out3_data, MC_kmpNext_out2_data, MC_kmpNext_out1_data}), 	
	.io_Empty_Valid({MC_kmpNext_out4_valid}), .io_Empty_Ready({MC_kmpNext_out4_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(32), .BB_COUNT(1), .LOAD_COUNT(5), .STORE_COUNT(1))MemCont_MC_pattern
		(.clk(MC_pattern_clk), .rst(MC_pattern_rst),
		.io_storeDataOut(pattern_dout0), .io_storeAddrOut(pattern_address0), .io_storeEnable(pattern_we0),
		.io_loadDataIn(pattern_din1), .io_loadAddrOut(pattern_address1), .io_loadEnable(pattern_ce1),
		.io_bbpValids({MC_pattern_in6_valid}), .io_bb_stCountArray({MC_pattern_in6_data}), .io_bbReadyToPrevs({MC_pattern_in6_ready}), .io_rdPortsPrev_ready({MC_pattern_in5_ready, MC_pattern_in4_ready, MC_pattern_in3_ready, MC_pattern_in2_ready, MC_pattern_in1_ready}), .io_rdPortsPrev_valid({MC_pattern_in5_valid, MC_pattern_in4_valid, MC_pattern_in3_valid, MC_pattern_in2_valid, MC_pattern_in1_valid}), .io_rdPortsPrev_bits({MC_pattern_in5_data, MC_pattern_in4_data, MC_pattern_in3_data, MC_pattern_in2_data, MC_pattern_in1_data}), 	
	.io_wrAddrPorts_ready({MC_pattern_in7_ready}), .io_wrAddrPorts_valid({MC_pattern_in7_valid}), .io_wrAddrPorts_bits({MC_pattern_in7_data}), 	
	.io_wrDataPorts_ready({MC_pattern_in8_ready}), .io_wrDataPorts_valid({MC_pattern_in8_valid}), .io_wrDataPorts_bits({MC_pattern_in8_data}), 	
	.io_rdPortsNext_ready({MC_pattern_out5_ready, MC_pattern_out4_ready, MC_pattern_out3_ready, MC_pattern_out2_ready, MC_pattern_out1_ready}), .io_rdPortsNext_valid({MC_pattern_out5_valid, MC_pattern_out4_valid, MC_pattern_out3_valid, MC_pattern_out2_valid, MC_pattern_out1_valid}), .io_rdPortsNext_bits({MC_pattern_out5_data, MC_pattern_out4_data, MC_pattern_out3_data, MC_pattern_out2_data, MC_pattern_out1_data}), 	
	.io_Empty_Valid({MC_pattern_out6_valid}), .io_Empty_Ready({MC_pattern_out6_ready}));

	MemCont #(.DATA_SIZE(32), .ADDRESS_SIZE(10), .BB_COUNT(1), .LOAD_COUNT(1), .STORE_COUNT(1))MemCont_MC_input
		(.clk(MC_input_clk), .rst(MC_input_rst),
		.io_storeDataOut(input_dout0), .io_storeAddrOut(input_address0), .io_storeEnable(input_we0),
		.io_loadDataIn(input_din1), .io_loadAddrOut(input_address1), .io_loadEnable(input_ce1),
		.io_bbpValids({MC_input_in2_valid}), .io_bb_stCountArray({MC_input_in2_data}), .io_bbReadyToPrevs({MC_input_in2_ready}), .io_rdPortsPrev_ready({MC_input_in1_ready}), .io_rdPortsPrev_valid({MC_input_in1_valid}), .io_rdPortsPrev_bits({MC_input_in1_data}), 	
	.io_wrAddrPorts_ready({MC_input_in3_ready}), .io_wrAddrPorts_valid({MC_input_in3_valid}), .io_wrAddrPorts_bits({MC_input_in3_data}), 	
	.io_wrDataPorts_ready({MC_input_in4_ready}), .io_wrDataPorts_valid({MC_input_in4_valid}), .io_wrDataPorts_bits({MC_input_in4_data}), 	
	.io_rdPortsNext_ready({MC_input_out1_ready}), .io_rdPortsNext_valid({MC_input_out1_valid}), .io_rdPortsNext_bits({MC_input_out1_data}), 	
	.io_Empty_Valid({MC_input_out2_valid}), .io_Empty_Ready({MC_input_out2_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_1
		(.clk(sink_1_clk), .rst(sink_1_rst),
		.data_in_bus({sink_1_in1_data}), .valid_in_bus({sink_1_in1_valid}), .ready_in_bus({sink_1_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_2
		(.clk(sink_2_clk), .rst(sink_2_rst),
		.data_in_bus({sink_2_in1_data}), .valid_in_bus({sink_2_in1_valid}), .ready_in_bus({sink_2_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_3
		(.clk(sink_3_clk), .rst(sink_3_rst),
		.data_in_bus({sink_3_in1_data}), .valid_in_bus({sink_3_in1_valid}), .ready_in_bus({sink_3_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_4
		(.clk(sink_4_clk), .rst(sink_4_rst),
		.data_in_bus({sink_4_in1_data}), .valid_in_bus({sink_4_in1_valid}), .ready_in_bus({sink_4_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(3))sink_node_sink_5
		(.clk(sink_5_clk), .rst(sink_5_rst),
		.data_in_bus({sink_5_in1_data}), .valid_in_bus({sink_5_in1_valid}), .ready_in_bus({sink_5_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_6
		(.clk(sink_6_clk), .rst(sink_6_rst),
		.data_in_bus({sink_6_in1_data}), .valid_in_bus({sink_6_in1_valid}), .ready_in_bus({sink_6_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_7
		(.clk(sink_7_clk), .rst(sink_7_rst),
		.data_in_bus({sink_7_in1_data}), .valid_in_bus({sink_7_in1_valid}), .ready_in_bus({sink_7_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_8
		(.clk(sink_8_clk), .rst(sink_8_rst),
		.data_in_bus({sink_8_in1_data}), .valid_in_bus({sink_8_in1_valid}), .ready_in_bus({sink_8_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(3))sink_node_sink_9
		(.clk(sink_9_clk), .rst(sink_9_rst),
		.data_in_bus({sink_9_in1_data}), .valid_in_bus({sink_9_in1_valid}), .ready_in_bus({sink_9_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_10
		(.clk(sink_10_clk), .rst(sink_10_rst),
		.data_in_bus({sink_10_in1_data}), .valid_in_bus({sink_10_in1_valid}), .ready_in_bus({sink_10_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(3))sink_node_sink_11
		(.clk(sink_11_clk), .rst(sink_11_rst),
		.data_in_bus({sink_11_in1_data}), .valid_in_bus({sink_11_in1_valid}), .ready_in_bus({sink_11_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_12
		(.clk(sink_12_clk), .rst(sink_12_rst),
		.data_in_bus({sink_12_in1_data}), .valid_in_bus({sink_12_in1_valid}), .ready_in_bus({sink_12_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_13
		(.clk(sink_13_clk), .rst(sink_13_rst),
		.data_in_bus({sink_13_in1_data}), .valid_in_bus({sink_13_in1_valid}), .ready_in_bus({sink_13_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_14
		(.clk(sink_14_clk), .rst(sink_14_rst),
		.data_in_bus({sink_14_in1_data}), .valid_in_bus({sink_14_in1_valid}), .ready_in_bus({sink_14_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_15
		(.clk(sink_15_clk), .rst(sink_15_rst),
		.data_in_bus({sink_15_in1_data}), .valid_in_bus({sink_15_in1_valid}), .ready_in_bus({sink_15_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_16
		(.clk(sink_16_clk), .rst(sink_16_rst),
		.data_in_bus({sink_16_in1_data}), .valid_in_bus({sink_16_in1_valid}), .ready_in_bus({sink_16_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_17
		(.clk(sink_17_clk), .rst(sink_17_rst),
		.data_in_bus({sink_17_in1_data}), .valid_in_bus({sink_17_in1_valid}), .ready_in_bus({sink_17_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(10))sink_node_sink_18
		(.clk(sink_18_clk), .rst(sink_18_rst),
		.data_in_bus({sink_18_in1_data}), .valid_in_bus({sink_18_in1_valid}), .ready_in_bus({sink_18_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_19
		(.clk(sink_19_clk), .rst(sink_19_rst),
		.data_in_bus({sink_19_in1_data}), .valid_in_bus({sink_19_in1_valid}), .ready_in_bus({sink_19_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_20
		(.clk(sink_20_clk), .rst(sink_20_rst),
		.data_in_bus({sink_20_in1_data}), .valid_in_bus({sink_20_in1_valid}), .ready_in_bus({sink_20_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_21
		(.clk(sink_21_clk), .rst(sink_21_rst),
		.data_in_bus({sink_21_in1_data}), .valid_in_bus({sink_21_in1_valid}), .ready_in_bus({sink_21_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(10))sink_node_sink_22
		(.clk(sink_22_clk), .rst(sink_22_rst),
		.data_in_bus({sink_22_in1_data}), .valid_in_bus({sink_22_in1_valid}), .ready_in_bus({sink_22_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_23
		(.clk(sink_23_clk), .rst(sink_23_rst),
		.data_in_bus({sink_23_in1_data}), .valid_in_bus({sink_23_in1_valid}), .ready_in_bus({sink_23_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_24
		(.clk(sink_24_clk), .rst(sink_24_rst),
		.data_in_bus({sink_24_in1_data}), .valid_in_bus({sink_24_in1_valid}), .ready_in_bus({sink_24_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(10))sink_node_sink_25
		(.clk(sink_25_clk), .rst(sink_25_rst),
		.data_in_bus({sink_25_in1_data}), .valid_in_bus({sink_25_in1_valid}), .ready_in_bus({sink_25_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(32))sink_node_sink_26
		(.clk(sink_26_clk), .rst(sink_26_rst),
		.data_in_bus({sink_26_in1_data}), .valid_in_bus({sink_26_in1_valid}), .ready_in_bus({sink_26_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(10))sink_node_sink_27
		(.clk(sink_27_clk), .rst(sink_27_rst),
		.data_in_bus({sink_27_in1_data}), .valid_in_bus({sink_27_in1_valid}), .ready_in_bus({sink_27_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_28
		(.clk(sink_28_clk), .rst(sink_28_rst),
		.data_in_bus({sink_28_in1_data}), .valid_in_bus({sink_28_in1_valid}), .ready_in_bus({sink_28_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_29
		(.clk(sink_29_clk), .rst(sink_29_rst),
		.data_in_bus({sink_29_in1_data}), .valid_in_bus({sink_29_in1_valid}), .ready_in_bus({sink_29_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_30
		(.clk(sink_30_clk), .rst(sink_30_rst),
		.data_in_bus({sink_30_in1_data}), .valid_in_bus({sink_30_in1_valid}), .ready_in_bus({sink_30_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_31
		(.clk(sink_31_clk), .rst(sink_31_rst),
		.data_in_bus({sink_31_in1_data}), .valid_in_bus({sink_31_in1_valid}), .ready_in_bus({sink_31_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_32
		(.clk(sink_32_clk), .rst(sink_32_rst),
		.data_in_bus({sink_32_in1_data}), .valid_in_bus({sink_32_in1_valid}), .ready_in_bus({sink_32_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_33
		(.clk(sink_33_clk), .rst(sink_33_rst),
		.data_in_bus({sink_33_in1_data}), .valid_in_bus({sink_33_in1_valid}), .ready_in_bus({sink_33_in1_ready}));

	sink_node #(.INPUTS(1), .OUTPUTS(0), .DATA_IN_SIZE(1))sink_node_sink_34
		(.clk(sink_34_clk), .rst(sink_34_rst),
		.data_in_bus({sink_34_in1_data}), .valid_in_bus({sink_34_in1_valid}), .ready_in_bus({sink_34_in1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_100
		(.clk(Buffer_100_clk), .rst(Buffer_100_rst),
		.data_in_bus({Buffer_100_in1_data}), .valid_in_bus({Buffer_100_in1_valid}), .ready_in_bus({Buffer_100_in1_ready}), 
		.data_out_bus({Buffer_100_out1_data}), .valid_out_bus({Buffer_100_out1_valid}), .ready_out_bus({Buffer_100_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_101
		(.clk(Buffer_101_clk), .rst(Buffer_101_rst),
		.data_in_bus({Buffer_101_in1_data}), .valid_in_bus({Buffer_101_in1_valid}), .ready_in_bus({Buffer_101_in1_ready}), 
		.data_out_bus({Buffer_101_out1_data}), .valid_out_bus({Buffer_101_out1_valid}), .ready_out_bus({Buffer_101_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_102
		(.clk(Buffer_102_clk), .rst(Buffer_102_rst),
		.data_in_bus({Buffer_102_in1_data}), .valid_in_bus({Buffer_102_in1_valid}), .ready_in_bus({Buffer_102_in1_ready}), 
		.data_out_bus({Buffer_102_out1_data}), .valid_out_bus({Buffer_102_out1_valid}), .ready_out_bus({Buffer_102_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_103
		(.clk(Buffer_103_clk), .rst(Buffer_103_rst),
		.data_in_bus({Buffer_103_in1_data}), .valid_in_bus({Buffer_103_in1_valid}), .ready_in_bus({Buffer_103_in1_ready}), 
		.data_out_bus({Buffer_103_out1_data}), .valid_out_bus({Buffer_103_out1_valid}), .ready_out_bus({Buffer_103_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_104
		(.clk(Buffer_104_clk), .rst(Buffer_104_rst),
		.data_in_bus({Buffer_104_in1_data}), .valid_in_bus({Buffer_104_in1_valid}), .ready_in_bus({Buffer_104_in1_ready}), 
		.data_out_bus({Buffer_104_out1_data}), .valid_out_bus({Buffer_104_out1_valid}), .ready_out_bus({Buffer_104_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_105
		(.clk(Buffer_105_clk), .rst(Buffer_105_rst),
		.data_in_bus({Buffer_105_in1_data}), .valid_in_bus({Buffer_105_in1_valid}), .ready_in_bus({Buffer_105_in1_ready}), 
		.data_out_bus({Buffer_105_out1_data}), .valid_out_bus({Buffer_105_out1_valid}), .ready_out_bus({Buffer_105_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_106
		(.clk(Buffer_106_clk), .rst(Buffer_106_rst),
		.data_in_bus({Buffer_106_in1_data}), .valid_in_bus({Buffer_106_in1_valid}), .ready_in_bus({Buffer_106_in1_ready}), 
		.data_out_bus({Buffer_106_out1_data}), .valid_out_bus({Buffer_106_out1_valid}), .ready_out_bus({Buffer_106_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_107
		(.clk(Buffer_107_clk), .rst(Buffer_107_rst),
		.data_in_bus({Buffer_107_in1_data}), .valid_in_bus({Buffer_107_in1_valid}), .ready_in_bus({Buffer_107_in1_ready}), 
		.data_out_bus({Buffer_107_out1_data}), .valid_out_bus({Buffer_107_out1_valid}), .ready_out_bus({Buffer_107_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_108
		(.clk(Buffer_108_clk), .rst(Buffer_108_rst),
		.data_in_bus({Buffer_108_in1_data}), .valid_in_bus({Buffer_108_in1_valid}), .ready_in_bus({Buffer_108_in1_ready}), 
		.data_out_bus({Buffer_108_out1_data}), .valid_out_bus({Buffer_108_out1_valid}), .ready_out_bus({Buffer_108_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_109
		(.clk(Buffer_109_clk), .rst(Buffer_109_rst),
		.data_in_bus({Buffer_109_in1_data}), .valid_in_bus({Buffer_109_in1_valid}), .ready_in_bus({Buffer_109_in1_ready}), 
		.data_out_bus({Buffer_109_out1_data}), .valid_out_bus({Buffer_109_out1_valid}), .ready_out_bus({Buffer_109_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_110
		(.clk(Buffer_110_clk), .rst(Buffer_110_rst),
		.data_in_bus({Buffer_110_in1_data}), .valid_in_bus({Buffer_110_in1_valid}), .ready_in_bus({Buffer_110_in1_ready}), 
		.data_out_bus({Buffer_110_out1_data}), .valid_out_bus({Buffer_110_out1_valid}), .ready_out_bus({Buffer_110_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_111
		(.clk(Buffer_111_clk), .rst(Buffer_111_rst),
		.data_in_bus({Buffer_111_in1_data}), .valid_in_bus({Buffer_111_in1_valid}), .ready_in_bus({Buffer_111_in1_ready}), 
		.data_out_bus({Buffer_111_out1_data}), .valid_out_bus({Buffer_111_out1_valid}), .ready_out_bus({Buffer_111_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_112
		(.clk(Buffer_112_clk), .rst(Buffer_112_rst),
		.data_in_bus({Buffer_112_in1_data}), .valid_in_bus({Buffer_112_in1_valid}), .ready_in_bus({Buffer_112_in1_ready}), 
		.data_out_bus({Buffer_112_out1_data}), .valid_out_bus({Buffer_112_out1_valid}), .ready_out_bus({Buffer_112_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_113
		(.clk(Buffer_113_clk), .rst(Buffer_113_rst),
		.data_in_bus({Buffer_113_in1_data}), .valid_in_bus({Buffer_113_in1_valid}), .ready_in_bus({Buffer_113_in1_ready}), 
		.data_out_bus({Buffer_113_out1_data}), .valid_out_bus({Buffer_113_out1_valid}), .ready_out_bus({Buffer_113_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_114
		(.clk(Buffer_114_clk), .rst(Buffer_114_rst),
		.data_in_bus({Buffer_114_in1_data}), .valid_in_bus({Buffer_114_in1_valid}), .ready_in_bus({Buffer_114_in1_ready}), 
		.data_out_bus({Buffer_114_out1_data}), .valid_out_bus({Buffer_114_out1_valid}), .ready_out_bus({Buffer_114_out1_ready}));

	elasticBuffer #(.INPUTS(1), .OUTPUTS(1), .DATA_IN_SIZE(32), .DATA_OUT_SIZE(32)) elasticBuffer_Buffer_115
		(.clk(Buffer_115_clk), .rst(Buffer_115_rst),
		.data_in_bus({Buffer_115_in1_data}), .valid_in_bus({Buffer_115_in1_valid}), .ready_in_bus({Buffer_115_in1_ready}), 
		.data_out_bus({Buffer_115_out1_data}), .valid_out_bus({Buffer_115_out1_valid}), .ready_out_bus({Buffer_115_out1_ready}));

endmodule

